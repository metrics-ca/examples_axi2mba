//----------------------------------------------------------------------
/**
 * @file vf_axi_mstr_mam_cbs.sv
 * @brief Defines VF AXI master memory allocation callback class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_MSTR_MAM_CBS_SV_
`define _VF_AXI_MSTR_MAM_CBS_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
MLdElfjenVX0yLRDL7eE70L9ACpvdxZjTHPyoT8E0qybSkukYxt5b5Q0xrDHZWtw
BSK5KDYYTy+PsoODxc25Wffrg/qfjja+NmDSAZ7EK2oVlfw6sCvKKK02b+6aI76w
v6PEEUH4UekJaawYi3PKDp74ZwM2k17Xbk+hDYA6JPsg4yRQX8JLexgrb+/eopT9
QmlZ3DLSFCY+kDGz0KuPqqxR1tGlIZ1b4r48HQQbelmpHX6HHyiCiJWgA7DY0NkB
lWYDLrp+chs3/YOOIOUpkvHnMstFJlJCA2Fs3cnNV9PEf6smSHGRxeldN+VVQNCF
VKIas+wu/OOs5cF4IUlS/A==
`pragma protect data_block
80dp9UdmZYT3cKliijcYLrUyQisAPA5eqrDx6zxtU8Imyb266k4xQmqLHBi9g6Lh
GAWvu2Fa6DNX+vKLDVhWoXf/IAPB+ULO+QrwzqXcpNAkSoPJY1qGocRRNrO8wUSj
7dQgw6vnJw7IE0zLfTU5dIxK+Uj2+wELfDfNyh21lJZHeAVla1NJlinE0gNLdcIu
jmQrgV7bpo5J8PQlkyC0HnS6aJHOjJTTz1m+YD06pAHJrNjiz585RV3gpKXVWxnZ
XTM5ElxlqrqHTGVDaDMaMcD04q5NCBBuanmeEfhih/CgXWF9wkUYMdM8alhygj8r
lKTmbiMbzoZIKG6h8XwRY7pEHLOwLnTlk0OUo86h7fnzF20TdHNZyBfMb9FqWkOk
q9QegJYHMf1jKt/WRgpHbbREXog+eUWJJ1qWypv+oFAxYPbRMR9jTByoDPCMd6pD
8ydAJ9iPmgMk2yKwo3kwRuA51U+kP3dtKDgFK9eGscz4fmDM/qzAe56a1u13omVb
te2rQydZm9m0pL3tWLW07856oQrcuQMKGUMGeMlwiu0v0J5P4kG4XLFkRVetz47s
zDxEkwma3Y6G0J16kAR4Wt7834PtunPpWybWo7NGRdoA7OSCtLaiTOv3sQIkW7m6
V7NXZ5H/G1IyNJTdenSlQ39bsfFRXCX4AAzsawAv3KkQIZZGbDh9cfoiknNMJe6V
V9KZkHyMpVFbTH+DpsPCAC0PETOh+sMpF0xTC3mu2TvNXl/fipK97zH72rHK9jx1
LazFm+Wa3iY7BYy+mB7+VudZD90tWo0A3QyKDkExWfp9H4eD7nVqPCF/8pS1Ua8B
DuCNYEqMswnFh3Df1qdPe3gcTTWal5Ug+I9eoqjp8gqRon7MXUykLcW6NeJWhfx8
tAEfwx9OJmUraKvkLod8yY5XsH5gGFfSxRUbLG9Vlk1kV+ACgr85NNwJuSXkpFGI
Rfg0o4/rBpAQzuAEkgsDsuAlykIjZgnYYlwDhjZrGygsMKfz+FbH+OFymvARDbbZ
JgHu0Dmsf3IK/QNkIokwcZODQ5+22R8AcQAmKZqqr6HsSSE61caFUBrV5YdUuZUA
QJ+ksQrTDp7bToRraBeNJdSTlzRaQmHHCFcumAipqcltC0FV1croW8sAOKfpaRGM
uc8CcyHCoKz3stE2ORT7Q1a3sdzF9DfVj2PgLvnIuUfIV0TsL+UYgf/Uu+WXCGCQ
MQm9ZwUIis/nkHkUuTIfRTh6HWcAQf+yL57Z5+yulUU2CyIjcA3+l7PgLVgqskyA
R6liX2GBSJvHzXbge9oWV3RN1x0EoJd8gnTw0exVAW2ZHCh5+f4LlAh+h5BYEbBD
s2Ll9PMGYkEhurKM2h/ZDYEfUpHmZrbc2JHXcKch6TnG7GwghObuIAXyDdHWioKQ
He3WRL9SxMSEkGbvvhc26i6Rp/qQTMOXOGhZ3Off9t/boXEk/433nSECL9T3Z+RK
vZR7lP3N6w4mKmWLFyVz85kFBD+S7ca3rCHBo6Ia++C3JRQUqiwKonTkwsqLpubb
9I10T+G5/79zzg//seFwwLDZV1g8HR2GRP08El6Ue7KLxPKZHMXTf74kwrwnAaEE
5O/y8LkwfhKIXIy1Cak4uAFnog3cBz9wZyVykYX2B6/DuHRgUq26zghQ8Hpvz9VY
rjgaUAyB+O/iKUNAp8tAn5w2pMxCxIk+yucHEzx3Z47fAr+EBmzspO5kZuCH8Q2l
xMwM5IdPwzN5yA2qSObhapaXLzB+lij0TNYFhG35yNVE6BngbcK4eVGV07rBKr+s
vHkNcbVe+WHEqf85dN9xCARaejOciMhAGNCRn54dkhF0ty01yx959kE+5P73qrm/
Ho+c8YAEpiaMdzOD6i570PHnPXr/vvbnz5tbmW7s2OTZ2oaJmUxCqi3KY2Q8uSXU
+a4e8vUtlPZ8d4h4t8XwhuQCUIy2A8hMaT8pPghAF9rvF2MUd+u5ROzF+gCb68Ia
m5InXnXntDEI0nYVcDkgqfiN3UnwNWVGcBtsb/3JN//uHuihscKZcQUdMM42Z3r4
aTkJBggXRu3XOBnOUDqgPqDYSrS5iGrdUZn5WGUzQuQgxfGt1Z5SE1toZE/mh19r
7RbbkL6bHOwz6l+u0jAYJZz7JCnnFiDet0y6BhYei25XKZWkLo/Xajd9G0XB62ct
gppDiguqZ+BTz6r6hQU53F2dnVAe2EQ/x0+oHhBQa8d1zKpdWKmLsJkXHariaFCD
oa6JbDs5mv3TXIq6pOqBY47A+onePkhymsl5T+lnpL3pD7K/IguYheV2CO0GYoH4
d6ZaF9czkNveIc2y9TfLPCFhYWF5VSe4m1BTN09kMLC6siTrrZNjPSZj/TFmWdAH
JMGv6pQmfWaPb8Uyv5/be2EUHcOrRH+dfoAR1Get846QqnGWUGOE07Kj5aUN1Ewj
4CNbby3EWixWL1MYenlaMSz+lRHeP2r2KCZPSLXBrRVYLU4z9kdVCKH2xFRRApu5
rqmtwSb0HZbvzN4XmnD+d8L5+AyY6bx/NkrZlmMw3qTEskc/GN8U7ldrfNnKg6UJ
ABT/zvJJ29tVbs+NE5Jd0adOHVVvfqrkna1xXfUJ+mOGadYKDX8cTZsXg1Y816Tk
GtReXQJMmyxI5mYBYVU5VeF7B1yVLCp5VJ8GUAG1qXOYFnmPgjp7KdaKp+RU7Q0x
l3hjG/hHDKveSgFr4EP1Iw6H33e7xnGn3SqOtlNe0jUSsPUElx/JIiRWMr78Midr
W0fxS3UtSm0CVo4fk1uTMbe63BPcqAig4CAb0N0Hu5bBPdHM4fHDnUcyCK8uWf5x
KgMJmoubFe36k0kYWcY2YEWrn/YC2YAsiuUu2VyxAkAdrZi2iXtCwSY7Z8V4WRuB
AmX312UMZ0EjA1QFI1UvT2J5X1m7By9cw6NXDZdHXDLes24vO8oL5Yf0JMAN1NO2
BCOr/Ko4a06GWnaoHQNY1RFmTOsNoAstlKo6d+M5Oq4xZwE1yFN5D1/CCqPzDj9u
yqi3bx9o3TB+qdz1usRp3GD8L6r8FPYLOOzTZ/TChBqCM9US4cu7U7pS42ASrcYs
FU13oidnzHrxQOPxD36/AhFhs+cYATt6LfXylkbt0GnHSbP9xAOTyrGoDLVoFGa4
H8k2Xz0vVDi3KRwrB2EzOv9u5bwCtAOkOVLNkZMWQEmkThUICOoAFGJtiO0DUybm
EfaE5cEwSEHafiWhaoOs/qyRgHLRHR8yJchnzH+fVMMVM0hN2iLNsBVpthBaE6U8
qxAXlaqYveOLWg7I3vEqQbd2YmQr3yaZdSAj7D2qxB41cMCosbUyh/WZmLIqbYrP
taTERsjUek6skJQNE9PNmn2a79GmbLRuWgrW7LTPbGQ2/3hx2UK+mdAJbgRbfP8M
t1/ZMmGMOlZNBUmTXDPUUL8Ou7D8IqRmfeWt9MssSIuPyv538eur2zLCAuBN+NyT
6RxBm7RwjWiiCJmKW6HZW302BUIN+7ghdMI50YAd86o6MysLQpDBZhPWkiuGDftB
jgDCfvsSTTndeQxXn9bqEgEUs0at+an907JmrfWgySTJ0nDbk3Oj+HM68brDIaHZ
z3fh1Lwi0KWPpHzJPdErVgtULUvJ4RGb4Sd8KJaU2mhktxNntQIvFllSI0JWR/nT
wM0tO4HKie75AQBhXQ58DGVtc1TSa156ZJOFue8NNC2YXubAh0ZmuKaP/M2X9LVd
iCz+Y10r9ggiPchYm1DJFe/qc0dvABeKcBMrDN81hvk5xZsXMrxBIntpjdb/f42h
5b4KIG2fsUiSiwHkLoVKXxi+zq8YiyzdBGjh3QHTrDxCIOdZlj3Mg94xicxFONXP
w1uSwThWnD4fkkVhKrv0K0ea6IFWPPAGr1dpDDiqLr7EHU8dA3KxyaW+nbJ7K6fa
IwBViaiTEDxIkO+T8cSed+7zgTt8CNukClLOgjQx6lcOJajydIOYZnlMIdKf+Fvd
qAd6LiF6q4hlKscLfOjG08Q79Vb4GTZC6ELF1rMqVClZ7KxZsCkJkhiE1nLZKlBe
fSQgdm2+qQpijnziJcpJn7C5QpFzOSChPWfuejSba+ft1z0Eezfg3LVlBgE9ZID+
2oGewD0fMyHf+fH/glFIkvGVWSWw8mCUbKyp6nRuDcGZriZAD18K+QXFYQh24zKH
SonOpRuxDp/ftKZ6aH6Xr8dokWNb2G3S7uKwVohtfTwdeVTliP3a8GHWPAciIe1b
NXlc36FwXX9uBXxBG2tJcQBA57QbAAfB4t5C3Ka3V1ker0j5pYj2s+zTzfepDmSp
W2qWAW979Q7nQYqavfKee+s/2WajNGM1SWa+hvUz9+8DkaeNXFamHVzhz2DU4SIc
nBqhDXQ8+CWOeXZdgBPNhAPKpWrL1ajW/WNk+vcfskCkmZXTqmzldZ0h7jr5vnOj
fJ9oW221S80Edht5cSLsbI+7RGTqMucvAfT2j01eEupQagPYizjhdCNhN+PkjiCt
AyTSgPuI9ncal4T3tpkIRZVth2YJV2aXZKvR3aDHQ8B2NwGOF2/+D9GtePdqCIl9
Pax0q+0ZqgykteiKqKzTlQhH31eMkWwORKyj+0Nd+TwI9b/Jmf+Mlih5pF2yrYeu
hJVk882orCHdyr7psS4HduIl8DpDel0+K0296RNhQo+7ouAOmY+HV+aYwTQ0fRAC
ri4Gr56sglUeZyu6LwdNMA+XOS78QKDCOI+qG5Qp81A+lwL+TLxzWm8Xg8jBWJog
7nVJ3d8oTrbv4U7dGZ0llh75pq9zHopELdwiqNyFguAx5CT/dUvJmy4Fm9fEOWCW
n8B90lMcvvB6Z0GrAfM9SOF11k/BV3PXGcD0wm7LlVQJFFW01mR94ccJieVou03C
4tFEj4g2x/jUopv84+Q+Rp4iJMNyauuIrvaIlPpUZm+RwKaFveJCvArVUgsPWc3a
AjIoBU5XjnnkVpfj8NusvVxNPhM9TfW1VgZKPWZO4RrdG79CdLoSmmp/JbkbO6IT
LLZ/GRJZA2GlvRaIdvWe8r1LJWzyMUxZfYDAFoeLDUVxXbyFAIU0nDiUgvMBLGoX
HzRnGPwAcqP3RYAMcgPJkcv4N088eQIzmg2G6SeyGsbvQ50vRAxcnS1WLklQXMui
lhfGBVKWBjwU+xjuqzB5L5yAm0nMSHzSsJK7/dnS1OyDJ162PXaQ1hrP9XhbX5Ay
rrjlVGMP2++27es05Of/5JRYJifcdkZ0xHcILMJytEZmru5rLtZfvSyyeuRgEWSs
hDS5JXItjI3OMkWkV+iORLv2xK/o7Rqfxm3yhKTGq44BodFZmzWLnJZQuxLT74xV
1P5U8ipWxUP3zGinPUrlIzL4gbo+wkKnVZHSwi4+gvLL8Vp4KoG9jXbiE5d5uC3W
ChkUfrAyRJLOmlky4G4ObmGRmeXr3LtCda4tmkcYTPBAVEtAQ8t7N9IVKbjr23W+
OvQLIxU8466rtgNEYD8UqndIZjPkVvpH7t/odD6niI8xfYW7B12falHJVLQZodmw
1EtTmKE7q6+lT6MXdhbZ6k4hq0aGiLr+b8oKk3os4SC0CUnzHWQ3gNJjx8UQIiPI
EPrwh4tyUrhOhqP3imHDHmNMFFm1UT+LTd4qPv2LEfGbJ4aaP2CR9Wku+uzvHm97
yuXkwpDiI0Tie1xTkghX3DKcF6FBsBtTYwnKI2NKuo6P0OoF4rt5Pmi4OtYUrPz1
ZzpRgT1eKlqm5wPxNUdqjxM7s0QdTFEewrIdGq1oO6CpwuTBzwYcQl/3IP1ZcXbR
kAvOAYsR7v5quOoRawulC/mJHumFWd1fNj11rGWSQA7xFAdpzf+og6WAZfMMAVDz
ZZTFM9T4OtqJDKiBdZRd+T9Ir9oXiZ+AUNVd1yELTj7OJWPtEgaQ88R8iG87bP+W
jNPssNKv4gJQwM8BNObb+1VDsAUXGrn+YzWH/O5U3qxykuMF79J5k4IByfgTTFO1
U8Bd7abvLsrDzmfLRzwMvZMjvZKWeeJN0xcq7jdVTRRCBNdMXvtdevYUE5gULJQp
c4+ileztmCWlg6l0u4Go+r45v6pG8GT/wb2636c2uEFQAWQu1ISYQMkby4PC8k+O
lfKlYT4xsU2bORAp+h6LWWRclFkNDUMn51phJ/SHfa3OzybYeQ57boEZVQG9pWPs
Fk2o+NJAQjWX8O4EhFVWWX+MP0dolZ0uM3obcsna67L/50DLacHJ91sEzLpkVfba
xLo+fhsm+Z6oOF4kjoKUQv+bCCHN0drZodhklnvOnQRGPHda6kQkGHhJxqNZxUkW
jMc4ry3VVb4PbJ4k4g5WM1QxDjPgjLwP0eonTt1FG8MtfcdZugm8fTbQU/w2b+Vw
2MS3Cfs1jMgb2GFw4hNC6zU4l0YEkaONoSLGnl3GB3AOAgdzkqHx2SQmG7kqJq4Z
bdBal+GwWkHxvWwPcA/Q8WW4Evjo1OhYFVxdw2yWPQY8/aF9MaZ21pGuY9f8TSIU
4M2gMcWcqmxrxVg82AXnDhs5ZLphIBa13rGgO1mvy60d4HL3lWf/A0O9vaAIRSVD
6rSRNnprrLHjvHM7tEELcAedm/cveU77qzCAXsioifYAF4TlZfT09rxTh/AbGTef
a1bt+V948nvkH3dHy0R/6xjzuBZkGWfYe/nzXvQdMsxBp5M7Rp4F0rCQC7eBxeA5
nfefHK+xXOK2/qbxgQ5NK0GqCTRagAZsrhxPt+/Ft+2wDB+0s0VxzZTqILOBDiQ6
+MOCv0EV/e8310Mxe1E9cHvGEy+aiqBJdlwx2daw+pI0PqYQSzNYLg5KkBn4QlRk
ScfIg5ts6oeySfOEuV7C9N5VFxDC512b6X4RYioyFO8lM2za/vBQVXT0FGRJU2Js
9gwev/yZivVaMEmpTUDgN47MqAdsED38RGLzWHe4zmcxjEI7ys1MxQFgcnQBrxVK
4wujcYuY0NuP6VrnG0U8dpntBFJOGZ4J5XDbEK3Ob5i1ukyUOA0VwStMDFK+kpbm
XYQDDMPZ7xpbPrJW0pYZN6gosVtvuBn+6NCzr9yzEwJeFmv0HfPSPA0vlUHi3rBx
oyvOOpcwKM72UOfTo///YUl9kV1jtsnp/zZQODKoN902lgNBMVxyqL9++CCFxwye
gbyRLznKM/JGlCamchZ12rnd4DcWz+cMyfN84mHovTtXAzNLlkAs07A6uVBPap1R
biy4I3yQVi2RoKBaH4D0JcwmX5Jd44/fnZhSv1YMfcOPnl0ls6cnqh85AHYAmtvb
31WDUVPem76sC7Dt/Mj5MAmDImVlGN4npLZ2XRyw98IAL8VylrcGant385RReii4
l3cJMCVogK+uea1sXcEyqECzjND1VPzddnINO0ljeyNMDl6/J6ezTNmYkRIKHCAH
`pragma protect end_protected

`endif // `ifndef _VF_AXI_MSTR_MAM_CBS_SV_


