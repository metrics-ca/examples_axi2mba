//----------------------------------------------------------------------
/**
 * @file vpr_q_typed.sv
 * @brief Defines VPR Queue typed class.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VPR_Q_TYPED_SV_
`define _VPR_Q_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
OBhdrK+XJbUY8PcN0+Xh3V/SsEDIA9QEFh4lgd2XM81SrXWLUxcLbEVWCOtFmQQL
k8Ufm4gfoYiJ2pLtfBYCtikNjjY8U0eN3ZWmg7BBC+JkKcFsVAz600yhp540VjZh
tHMXhJfGqcvSvPYfLq9Rjabd+7pVHJWE3GMQ+NFiR2G+Ge88ESnTO4aq0VGU9QZi
upCHebViGUNR6ZZUzFIZQt3pJXFen7TRP+ArsALE/hc4uE6YdufhaAucV2wstZBf
Er4qexafVPX/FVUfqdEkQXHoI0gO0zHvdh3Zwh6hPC643Putozdj+iS0Fa0h4Ouj
bvn+wMdtQLmsfEAA6a7u1w==
`pragma protect data_block
ChQFFME4ZfoCRqPxBuRXbMhryZKFV26/WuIWWx5gh9VN7tmvow/zUVwlanVc2Mdk
Qsw5GcyQJS7ol98E9Nnn1zzy2XAid/5UvXf7GL1pacXl1aqSsYsaxP6DUBKFhmDi
cmCxI2MOsyP24ErrMY+mommTXFLznXHsI800W0bMAOILqdu60Zs2BBWTDvHEIxUP
Hy+X5N/pOUgqkCxZn/u0xZAyJVkqtKFMI5/d26lp+WdWkoWnm49cgEbsZxctormR
DUzrL1xi7kfCh2TADsF4gaNOceIxrCxuqAWsqZ8eLUmY9s8u8loxog7rITqacTtO
wYQTKo2Kmvo6l/nCo8l7P0biewYrwazZQUdYuvFAMeesEThrweSFmb4IKatNKPm1
1fxZka52tUoH94rxhCkLqoWQwRg2gwi31tcN5KX6EtgsVyAyu9RBcdtW3qCW95tR
8lzOSGj2HM9lAxIG3OEMSdQQyHXY7GF04EHq4YWj+MIZ0tRCCSVyIkUSg02+ivYi
/fjw/1+fH8K84KjiTh4GxNJo/o7JhDkodDGOvO95+FKNMDfnN72IAaV8ExkliGk9
OAZfVY3dBkQBwMBS4NjxrOnPNq3zS9bXxl9AESj1EsrNgW+IC8IN8hvaBenHP3yU
rgc0slVw8W430i1/yPD1il/vq863kf1qtrIYNf0a4v6FMVOcgP8LKDwb6Hv31emY
OXsNrLPTOjEuV6CtE55InR0Q2dBcgE/hR3MX/XDD3edR0SavPNq265jras069Rp2
bUJTwS9Fdq2Ee1PEmanV8GV8P2SrHitgG9RU+iI2lF7Uy8FOvsQiL/XqKLj4A/gu
nQCGb1KOCIp1Lrd0H9lqovXMSdwDxlePIkYn9iqrAtyK8e/FGSfOj8DgzDOLxvOm
xAed92xomIGhzXLy3cKNajWq8PxQwrqUwql8CE6qEcpgGJQ8zJnatUf8tZeKn4jB
2W9ElLe2iKtR/5ak6LoyFlWuw/qjglO946It+RvdO6RjGGL2NxWnW8bPqFiAqFyQ
NrgXfOG6cs+1+ZVNFh/TBEjwsgVpmP4skTznNFTMqZ0893VWRSOU7UXMeuyFLkx3
allsqotT1zE6LGVOCmKd8vxq4FyQny1DQkCBHkLtcmG1F0N4qyretPR/TBEGBXhu
ziPmeRy4hpl0sIt6cQb/G09Jxgy9yPad+iQksxea177P8bhq1lU/fzOHXqL/560a
hf/nc6h5z849+NyTV8zC7YCIIf+YwYryYZnYCdjXTiWf7nCnkhOFj76icDT0lyen
ONoZdiNLfri6n538tmHNA3CN56fsY/aITtIUy5+vXsbo5lApHuJbBFgXNbR334mA
AcyCAC5F5mCHdI/f/i6oLOZOxLZh5VESCCcZrI/BRd24MTGUdisD5ys0jcxhjeEC
gr8S38O4vxYxT31jARreHFypAy+jSdVrpXSlG9GoAkLLtlm/e7HPwBkSUA3s/Sfn
UeyFQot1LEgEKseIq17iSAEjCKSrjgByeiRTlVsJTiawNibX0sUN5DQLNEf9Tt/N
zKAkGgT6Q4S14u+hbMcJ8s8S9rYquCuYrhGlWCUp4xsNTuYzixaXQNGvKDeDPQKu
ZfCcLSpPBYPUX+Oag8Z9drXOuwv22ahVTVvL9o7W363OnMJEtBkPM6GCLuwsrKyz
kKPlO5b+0C1u6L1GJ9c9W5Qm35B+TwuU+/0zKs0B3cj2LSuJ5iwjkwIDbvMDue8w
8mx6QxCDQ80k7mxnq6iPzhl9dCShhz957l5lj1kuLPb/bGdjkGZvVsW2AZv9QXdE
m3RsIc1plqHu5IzSBQVQ8d5APRu+K0n9gsJnrb7gA+HAkCfS1NpitmfBhOtYEEGa
jrM52gDN7t8TRPO/txQQV7mqDrHD/7L/LCkGbeWtdBJJY5Wx4PD7l/q146265nKn
kXx2ukgiaUxOW+XQNHaCz5GWPJD8P+X3yEzIW4l5mwfuDbGK62W3NYc3GlGpbrHj
9pM4sbjJcqj4DgYV2oQHRNreO9Hux4siz2Y9PWGkbwr9My2cA9ObVyipKj9F1Awn
VWK22Qn9uHox7vw/rGeGxAF/MDgpiM9Blp9UVW68hQwZ7g2LiyOM5SYuw481VMuy
mPnl5M/bYP5ACRakGqyo39Ruir+WfjHV+LzwnERV0DKIul8levc8sZMrZF76pEP8
kGPMijqPUqbsKul36AywOCIFH4HBVsjsUDedpcJE1DOogny3NtRaRISon24x9sts
fOnqi6R6XOTJceSV+cDjW8Y2O5gDbajcnReYt+X3s1BfmUCFYq9bB5lKV8m4cwH4
TtX2oOzJN7QiqthLhdxyKsitvAGoVAUBw6U+bYPZUBu3xkMaucX1maIZsSAgYD7F
T4bZ7qsHVFeFNhhDUohn8KLmdQV6cgILRmJs0cs7MAUA47u4+RF8flqhzmN8OHc/
4lMOQi1qM9BxXuBRiMGVe5/Zyr5NCSoJdUKZdqGyAwMGj5amefYb7WiEVkpwKowB
WmiSX7Au9EdpPVMsejsbYErRvwH2UKpWZPE5lxwBKtaiOoHZ60SniI+/QiTtswZb
BOt8GwRnXvqpRxpQ3PBPCL+VBHlx8yvMcjR0nUIzElvMJjnD8POLeoxKz7zkGJZd
a4LBRoErTK4qX/uP6CJ2MU2DgW69Qkcy9M7w29I4lI0dGY5lz5YrqNFBit+cUJLm
FQCJYLIb9LIA1VWu7Lj3dS9wy0PYrFccFE7jfpMIBRRMrFFSl5gUFh+T4CCxnbrS
zPvj3M0pLohfpoiITrPWxPM9H3hQikhANvkYqf5MC6/yPohD+bNUSG6S7YUzOmb7
9mhxd7/MTqUG6Q6ga+dEWi9kHJuhfAvSVZZCD5dToIdbg/ppT60DbWolmhMPytwj
3ao9WC+ECrOsDkHqRrydfzmIFB6rL0ggja55etUUeGxgDk0MNaoSKWNqeEaKfLhz
LFzA/NHLCBZPBXw3/+uiPT4XLyCa+bGUssNz0TiLeXRyaZ8fZk1KZe5y6D8Wcobc
mZfnWjDhJwF4dntc7VNxkhZ4VlzpJH8vxjRkQ+buEh8R0UhKtiDktgJeHAhIVvR7
VsJYwOdCCo8BtI62E5EppQVzvp8Aip6gTUEFbdOdBOD503mKI9FkvE+yCRHHl/iW
wpEb/zXSbgl0EeR1U9WnOD0OFVllPre9Fh8cWdW0M8WkSgOOqCKrOix2EwPjLRAH
LlV5Z8ndt22Wb81Fmj1cjngqD3Go1oCVJBzV3/lWoO4ZN02cPKc9Ofz5o32wis/J
rH63FBqTpJA+/wsiOQbKjdcwyXD2Njr+x4vev0EEvlU9Fp5nXc+d5QbZSUua0EV5
6W4OGjZDLNudlR+Jm3OL/Ib2AhIK97YvKXQ59GiG9F77s/j4ihpQqFhhdEZnR+RY
nBISqyiy+S2iRX/gCNSX7aE7YDGyOhBEDWqsn1m87xhnHk1H3SozvFtPAuw9zBLK
bbXKQWfoyIJAq1t2ULNvBtSs0x1UqbUG0L01MpzikZums+wJSvlPLLPUI2lAgIBy
FO+2JU3SrxQv5k1lTz+BEHm+j4bOb9tvw9C2PL9F3UiG3nHciD+5USLjYhI1g0m8
XVK7v6YSXkLe/daiB9b1YJZXhFtMQZ8Wz5Y939pCvNCP8shg2oiA0leL0h8ajxrU
oRTey6e6i9XJbfo+qYS1phjPPIfhLTketZA9iA/xxURpvdXJJGJZblevDNY4+g2e
oeU9HyhAZSWerHlNhXqORPe9MWM/IZw+ql1qGkyB625JcVItol8HdS8Euww+jVEI
OBR5wKneDByxiup4cbePhJ2TeKtKID2YTjiz6xLBVcKbkYcMrWnqFHpEX23feT8m
+PKmX1GJOccdyoq1SCRNhv5p65I33oQ601Va6GkDMKfFAZQzdZSjVKj9cdW+7+WE
+8VwVW+j0aqQl00PMcHhUqYzCJYD57GDs9o34EZe4nHKwknLmlz0vj8rCacoD7Tl
8jtjrJvyNSrCtxhtMtQcBC3D7y7Coa3bOM9eb4vyHHMc10t4rZUUfqAXpXto6BVy
jJdPopX5Jp92cBPIY5JZWHRf5hlNNsJW7BVjo4P82Cc9HuLss63JNVbQdN2lctrT
EM3JUz1yf1k15Ojc/BGHkB+9PvHZJPkwus1uTDXxibHiPDOaMFOCI7cMDgsTDh8q
s3/7WmXlA5mwjbp/Y7Ugb0LenD6RTBTD2dEId5tOIVb8vutgERPtXCZwNpQNv90a
S/1iahQu0JOzn/qCMQZCmtwrKbYx/p0jvkDO2DgcIMU7WerksQ5lLebJE1uSYKiu
c60FuItcvLTFxwxMy9IhnSsVvchqrkflFKMPhyIz9/cAU4+/gr9ito3PpzEdf/ik
HuX5rPezithoweM+3QNzVcvHEJO1qrDdQPGeYeqXu0aV/o/YXy7Lq/TPyNOYCbRx
1O+OFTE2jpKTV86FIsIHgMN4pWEuoJGaVfhSzuJe0iWrww+UxM5R5mQ3pc3J+Elk
vncOwuCJzkVrofe5HPCs3leG7ngFsrf3Bo/CwgZfiBgQTJ+gYGkNms2mZ7vIVblm
7SJSJjPjhfbCZlru2CxYVjw+P8xAYQGaN2/b75ff+NT1cvJoSNTiMOWlUB0A36hE
VLNGCltD4i6Okuqz8mWW6Dw20qLcmxWKe4JXMqryqy2ruLzQHM83QP++oKX7Cju9
FnXf2Z2aHjJQLBfugmgtXeCQT3pyH9H9RysnqTNcnFdD4kcsQPgrxszeCwiQqOPZ
o8KI3wx+Ki5QdQYj1tuOcg3Yp8RqyQbm/VNe1+CSISsIAfdwXCEDKq1qWcCeeZl4
b70wzMlYHlP6k4vn4e4czWVklpjljSFeWUwf5EuHBzxLEhg5VWyiFtwFLZA4fCM3
vYTftbHoPRuzrsShWzl1olIryymeb3Yw9e3hTZEMwsTfNbrxPOmChTTpB1YuaEw2
esORSrKfPTEtMCW10eTBVAvrlErDQSw9A9DVvOQEYWOfhdI3nvgG6sf4cd5g3iRm
RfGlXIS7tdXGyc8zPhPdvaYV68qfE3pWyOWFA8OPbOLlgYXxoGn7YCqse5Ap7e2n
l+ZhgVGoc7uIFuTR1xjFnLGPQblRFJwRiyLHPUKfnkfEFnAB4dUU83Wb+gFsPbgZ
SleE57In34gXiWBU1wJjFBBjKPwjIsVdJuigiMSm+MBA2mJ3K0j6YXkE7pVZTjXx
ldM0CL7GKre8ioweWTd0IzIyAPTd2RCwtWg5TgGz8tIIFD/Yink/Jlk7f6DNo26h
ABw0aefhdIliY1ONqbZfNCyEHuMhhZIOCs8832Nw2cbnWH3HadMUtTsHzVYwANsR
nasJ5FisInpCoRpGEqP2FmmaTs9MVyVQGrMlWfMVhEXcCFm+uCVonF7C149hfWEw
AM+KQ23gId6TkLpjzmzrCCy4L229uQ0ikWF9HEgwMHugCq8RDJGRd19lyg1jvX/r
yEHKz7ztBs+p2HhNVPGRzt5/Lvfb4PnOIxCEakZ46tHL+mI9fdeHj0TuZdqvJF8+
tehTDQbvI+1vPcaDkzsFNXxokBFDuqOgvGw3r6TLxBsLNpAICXNWfb4VEgvqcBV8
9JHi/x3eazv/hBdDkPj3EtiRZ3xo6DQtOfiD5c6cCr43x18xBc6vbi7ajUb2JkYE
+fp8ePTXOGO5j/hjvpf1AJvP3cDkzntXMLsw0F44QcHgWI0KidzIMN1hULezMpbr
nmUyzvzDfQ05stWb07w7ObGE/9DEP5MA6qQovQpZ/92cGl+zVdY4+gESslZWLkrM
zF5iFWPnv8e6AmMqI+2BkZ84Y0voTezaXibZejup8IrOK0IL0dCqf+qxrodSVjhR
UkAq6I4arcIWtrV3G+aAZ1gNS040hBfAOJLxMUCMnk9LzoeUByYGY46pvnEeHn9O
xxBbZHJdvttyWqKdO5nV0HSgsfjktFeWReWuQvNg1+4xil7T/+jIpBDuHg9uI+8E
ap45LkdeOpOVzRfz/2UDV1M1g5j1MCa4cAg2L+4SvaW9/LJLqxMNEJZ8DirXx8Z8
RvSr3B24HcvSm/yRAE6qfzwy3zL6uFZlakTGATLoEb3tcWSiz6p8W5B+LawXdHf2
bAOujQ1KFOdrlI41Odi7ExeyPIFySjfsG/oHNvQWYpONLpk7pytoUf/ZAOfmpg9W
Ghbzib9TOwuzLitUDPSI8hKJ0iSdqTU8L4YKKahsu/r2r5Hu9lRS3dIBvSK6yCTi
A5BYGE+0bPQX/N2UvLkwiQ4zppqMxeIRvK0zLs02nWUQVKcgQeWwxItysm6UQQJm
FTkFEVwyMLQgnAwXSSGM+cJTFThnmabeA36jokt+w72ZoFmeA4rLQbvVr27DfGdR
8G284XmSyNORXYoi+J0WZn+ZHYJp2nPpClL3oPFEOQVqeAKLZhDRiL1kMjnaVZII
GcUGMiNiqXNToXp9nLDD/frfCeeIQzv5JkkVNo3kTeQXtuKT775sY+EccnLHxEbP
Z1XQLMnovb/qNnP+V1FrmQxtuDxxFgDEzbJ7lCIKE+HXzzEt0DzLQCygOq18KcKf
QV6Glj/K9GpkLrafz2F8gROKzPfW/03/+8datm8cC2k=
`pragma protect end_protected

`endif // `ifndef _VPR_Q_TYPED_SV_


