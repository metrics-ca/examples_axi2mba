//----------------------------------------------------------------------
/**
 * @file vsl_sbe_typed.sv
 * @brief Defines VSL scoreboard entry typed class.
 *
 * This file contains the following VSL scoreboard entry related classes.
 * - VSL scoreboard entry typed class
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_SBE_TYPED_SV_
`define _VSL_SBE_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
iAXdndu8ZlHqDL8ox07VNDyfnrEMZHCXHe3CRLnkReDWzauSyIuYJtz3T5V6Xx3/
koTiyARsPa0SbbTLT1m0yZgGQcyKrHvxKUU7pKJ5Zd2HE5kg82KONKPwkL58zaMV
yhMD4YTU+ZLlvGJp6iqipvLSo+UNfRac8YPGXukTHxCt6MlQuUEnLaR2aSjZqajn
yCTvQTZv5pkqABAeqs6fJ7Pn1jH5NuHtO63uFidO6TbG71MlzsPvB15dXFGtcEWp
SkAsx6dmt4DTWnpBWTfcmm2mpZGFzM8AHs0LdQg6MnTBVuQNe31aZ4y0hpUzzG3k
lWxR96Zbej8JYlJ8YsYLqg==
`pragma protect data_block
3STSht+91hWLwTzYbtLiZKUMCL1LET96+gvxfe0BMhAb7iQhRSvlzTCP5ZaIR7n2
SDk9sVPC/3GkonvzwsVfu98LYDZHqEnoJLwxyHupRi4s8epDSoNYQ6mGTU4r2YKr
JGVQNlHlrHL575HapGcRXgn816C1IDJm9eSN+oZ+08W7///6Wo/ge6LC2NexYFYV
g27NtljwhLtVMjUAsfi98eDId2kxyDm8e4SqpeCPG2Vc7v7ji9W2XltTQ1IsZXaz
/4jHv918RSo+fPtBfZPzdJVks9LW8U5FSnUr+wPnEspN1xwb0QGr16P5d69b8RdA
HBDDvTvqyFuy2IOYnISl4TljyK65ubNoqF4OplTxwXyDrjfq6GGONdV347vgM2oR
77zdkK6rMLr6JPqwjxQpWyQ83R1NpHj4M6BfkYgXOoELoJjbkav3GEk4YHHea3r7
TfYnPMzRAf3GcqxIKp9Nf5/npioQhdTXU9u+S2HLv+VUpVnxryNRSGkBcVDCKxv0
jsypWY5tPBZxaeXrRurV73JHvue6CI92Hk+lb9ERzAPTCJUQHv/JMn5SFXFkHFMQ
pnEp6vYPV/oERhDHNyA8T8Nux8nK9NGQY7WbR50DKFDEHUiMJSFZjNVOcjTsFwO8
uxAs/sYu+Z+mVe0lnTND9l9n9XskLISn9KNoizD/RepKkpGow4lAtaoKNoTA9fdM
QBt4qKpsqxNeynxE3bwYFli/A0ou8hy0wJ0ZH9nQ3tYAtM/9rbeYSWJVuAXMBavw
7+Q6BBd3gBx/T0krq/6nxiVM4msiu1fO5+rboudy/0qTFAh95WA6u5YNIAKWiqZ2
Ow0lOLSzYJwA2K6m1/Jr/FuYwkx2clxBjzzHQDghbToZipEphq12UFNXFAhp2bRb
yx2h/ZW+eEp8VDL8SOxETDOvpxzmIv8e2Kg6CtBUGkPZvwVt/uCj4toDUkp8sDuF
joZgTqsPWMGFJgCz7HkukIRgurKa8DdkGENUBSjVMrzEaz8BqR8++Gxv6Ne28vfB
NjM+ioHXQS46sUgIUco7ZSNr+iY3/uWCUTejGIlXgtCF18FUCsbvxhJVM3DBFXDV
moNDPMcwaCDanrH6N+RYcrE6XFzbwUPY+E7jk2EuOwYZ14YwHZrCZLiJehEHzAn3
Xka2YvlsIPaz+0J/PoA9BScqzyuahWpqT8Pec4X9z/ysDQKVB1Ltf4DKKdCl0c0N
aunChMX/y9p/WHCV/kclQ1BUIJeDZdHTc5cp3rYkaWu03dKS1GpQMwTYgI3lLCbN
hA7kyrT00bSycdPEvaBGI7W3Z0CCkEZyMTeh6pNVozDCnZvXbN+NktfgGZlVngL7
6bB/AUOcZiATD6cn2XgJGB96DThx17KdSufyBnX2WsEQNs+pJlYFg7ebwlMcJizJ
ybD0QZh27mtBA330JMhiMwQEoQMj1iahoTK7j9Ekm592CyaWBJHUJvmtBQOivLNG
Y7PIqxbyrau35n+VonZP4y4a1eK8Q0ZWhi44ntqXT8VjSTx7Rn1Lrl4EvIl0CPeu
SqQXxDcMMKVpswVVTe2ceh46FwwuBGBQH6Ng17sIU4Vzy1Y17P6Cx5H0MiC3ZKIA
InihZ8eJpZhSwXqinLW0gw3Q9IvWnpc0S1+yQ3/zgTIMcP0PZIRcEBUlva2NmzDs
EPdtslQ3xP1GdME5q9KS/097OeKXAG/6L2kS86xh9YweM5Vio6zm95WBkagIv+RQ
/BxNRbYvjNGPUpUkOruY9+yocJc8sB3bNZ3ASpsgGViypnx+KgTQ3k0LbwbDHEKe
PmlMkkoArbO4Xv+sXoHh4YKT9B4BA4mDiW7zyq0IW7LZ8rzmHvUgANvenDYCm1hz
92pNMM+Rv7g0aTj7pdbYDj5GinSLuW247JDCZVPoc0bddpKYnjzqTSK0UAO4CSc4
RdtYoRsQ2qbAfDZFbCSYMUigA1gH9Sf262bZtDCXiundgJoLTbfkrn34x8cq3vu7
OfbZWYYUu/VUyQzznPjHkFJV7X1xHn1YzJJMAWmNk13vMuTKDAJFyvZvw9Ny8KT/
aJa8lYfLltOZW6OGbuS9iBoAVDlmufCnsNyxuwnLM8GAVK0FLK5f46TXsQYQIQSw
S3NMG0b3skY1MlAm5nUfI/kiD89nufsUlg8FpoRtGK+cgXOqX6wmVCZZF+TCcgQ/
G3gSsL8jtd9dyav+3WbFUebJ2ulX7cyJqFbxSzBJlu4JnU3wb1HuhF8b4jk9ptXH
hJSGJUvmDwWLN/uUQKIPltvOR8IZQsdStGb7WKFK54m8V/T9MO/N27KARAHFSMKl
jPb1uhgeuacFpxJ9zvSiEpzfzsrDUcj/exXt6ROryT1HpxfHxiRWCmS36FbNtcbg
wccApaTFi4gZGjipX+OwZnJq27Ds52auLvPBxOSWbzmg00Bf4JVnH+7Ac/c04BXq
wICpXg8bnXpaSFG7oN1RlXmlvY9PjX3cZIh111iwkHJHCY8/LTqUj9yagZk2x3Gk
NhHXy/OJ8ZYVWqPLvSubPwcJ94sF68lUINl2BGSQYOIZqWHt2z9p1t69kdbiGiuX
0lJUoFvidqvbHMFE0b5z9ZqBGEuc9CcVdQbKpKBvJHnx0EjfMdFrrDBGX+OKHFIJ
ZNhuSMBCvMxx6mDult1XctC/REEuh6mS3+LYzfzL0eH8WKj7sfr+nIaQxF4p0FSU
/blsIufESgyQ6RtH7b/VNkfJTcaMawCbITBV6vtEwc2X+Dvmlzfxpw/2Y1JJBVHz
dy+lUi49nVCpZd2bBY2grtMGk0Hl8Lw+mom+Nr8/rILNHBuUzL2/QStQOC4LRzf4
+tEiBxV2QQTvrcu6287BNTcHptUfM+2s+wuXuFiPEm7hYkJEgStnreJPlrxsPjie
HByvpwCjayv1B2nhcd+d46Wu1QSqwde/99XeaiwkJPlUuiCoWWVYONS/6MXsv9mi
lahBU9B49g2IZ49L1t2th7OvTrc7tTXl85DJIW/n6H9tUButaJruulbJUzsAazta
lPQPbg/ousowU0oMAM5QfA88MDqQ9PCeBkaFtDqJnty+Esg1E22HQeR694XVaM6T
fxMWYgu9Aiq98fUjQo35oyY4B0r4ib9lVaaiU7iLzVndNz/vnqdBq7eQ6cEo7na1
eRAADZB0EIZ/ggu4gfmXeEpZMZ+/AIKGsmLP8PC98tnugF72Hk3kNZ5HkydfdbNQ
iTjmi9StsTHF9UpeoeB0wZ+Wz8dM7qMKMYWVuP6dLT8F0+kkgZnSp+uSA55UCsie
o/ccAXKjRRCM7O4MUblbGhHG3Q/QGR/5WdOrPJtGbxrLy7BCR2j9y8t+pH0j0sSU
CtKzCvr349PmbnhWtrABIjv+owojAErqanrUVcu8zKex9qy21F//Cm5bxeuokcQl
AR1bvpIY88QHzJDao8vF6gjZuwEDfKzJLkYpChDomaNpdjb05UY/32+v446AGz/i
Q1eJ0+FCH0KZOnJDSM/0TbZst6oQTCqJsEf67yOtrYp7B5ealYRVpJCZlg6gUChB
i9CKG6kD0TD2WN1IEAQEyuRGsAzGW0MiAPcPWGtVA1NH/HJ0BZi4DLzf3/LwsH3n
HcdxCJXZJCd/5qDGAU9UEMFvXnRSd4FbYGNrGVEj5OrGKdlS5yTjEiriOSXUap1n
NduePmDC5p0nXYBoObtOg12V24V/ILOLRftrgZmoJsRNdOIRCWAxrm7HW+2Y8VaS
1p2Ns8psfbUmCdvFoORJsKTnPSdbV1sMdZzTYtLV1BtW4CWw4FAhTOisxHoLoIRo
Wj8gcj7Z476b+iZ87IGM0wCrnbM/omY4VdzF8lxEAQRyHUDUdxSKiOPQceNdew9O
Bt+bxPQA0QDmfrqOemi+JXJwnWeckT0Qf0OVt7PTyGOSsxSbyLKMF+29EShH9PFB
ye0czc2OUZOE+tsFdQhP/KPbfBxPmGwFK7XvmNQ7475YtiDtU1+2tcsA+s2tF+Lw
eUx+gkH9fiQ0Q/ycBzpntNUlgYw5bZsQ5q3cGtk5COzqqm8ZSqf2dGzDWDYHzxTO
UcsiCHJISqSrIAzQ+XFknIdr0M9wElrgpsSfqzvXgs1IauARBGUMwm0/gMtfyZqo
GaaQHYMg3eru7dX9uw41I3etIx/oFrvNvzKFrp2qVe4O+9dNEg3/dPMS9lj+mV8D
VYJpYH1ZFeQLQhushuXuNQsguutpzypt1pEkFiQp4YgZmFYmCR/i7CkGASo/na+/
BUSv8EtBdIltAVUIUes9NbMxUqK0RwmF6ndbR6vDdpQ53V4Iv2XwwCW09xR7aSqw
Z1he7+35P5AASNiEsw8OHbpAhd/pZrhBb1MNCKq+2t1scNAXqALi2PGlGwa/c0jv
8+R6gDzeJhxn1wkhtmZXp5RTk7o//g0E89jM6gqtIEZeKYDVm2Fv1fzxPNG3FiCI
YGEK1k9eSD46fbGnE3mdzIM4xvWE8CccpXYwOnYncXMiAymvWFKkfevZYpqn3sxd
3IY6oqwKBL7EhL4Ml87QYtl3Gv2Uq/wDLwiMALBgfHFpaOBtFBr/caCoMFuj5JRd
zdGMp4F2JnljQKUqfLbv9eixX4bMYLpLq+sTfY+c17kLysQiMXjxFLNwpUDujFqd
N2nj+P8ES8gSXI7oTfEw+MOZkdfG5D7VTOUmcQo39fsc1A+exwGG8Kf6G3UbGfi7
qxg8T5gAm7NLWo8ZKLGRodiguYcODDTEyQo3p4Uz9UB6rMhbN8Ckw6eNu5/My1Tr
Sv0YUQHpW3EvpZbDMTkD+02x5HacXzYR9iql/NBkY9TP++ixfIzkD9UuxqqEEYHU
euen/hfj8hiZSGexnVkevTELdSOZHxM4FGvJ5gFk7veJp2fiGULPbWkZzyA9HJ7T
biL2/S8EbrU3E+MpoxXQJaO7/eJC1xYwl7GC5E3/hQYrQWIxJAbkVSgb210fWUu/
4c/mUgBGHsBScMe6gs4hGFuFRytA5YlS/+hLI2JzxlBu3l/psA3jOPdBK8ME5lAz
9RPuLDDQqAXNX/GomYa3hCGdSF+5yn/rzjfgN3P79DuZpXw5iqAM1ueTS2au/cz3
iRsZalkW49Gd0bmcEAZFlzLaGgiqJx7iwI4PWobnIv9m8Enr4z/fZmoCWBXdqLDj
qKMoiyp0ibol+yECSU/JKmPsfmqGq8Tc3qW3aqsR2BkK4/qNNNd5zXIVk75YqJE/
w6066J8hnICEOonuwIHCQ5cRpJvb93jsXsxN+cbbdu8/6QHWMarLPxKtOrKXFYXb
lEotoBmAmgdSFI5Pl+arwEbvwMBUnXcNhBGfDOed3ngD9pw5wJjPtRjRE8HwnxO8
P144rHDIx/HxlyzNE39N4J5WQxCW51hoNY1B8pUkGX/UtSE3Q6a5hWtBAkJEUbKm
qSeiXIN1tnv4pL3xdUxMJeQlZqyAOTpgOmc8lK739KsswGMCzc79ad+S538FhEtC
R/WfO4f9g2R3j/3X6sz/lfKvnZdRbQF+ZPLgV2noLFLTDrBCNaZcJ8iKUjUHZHAx
TtwNpk0h6+SZIKrd77OraHgWBL1dP3MrMgPCwj+yPz29LRQZpzwW4Xh4nFkAcGdX
A7HLtYoEnBW7gNvM7PbD+xNZSItGPYK3k87LAfZuR+p4F/Ssl1MgCvPqr3+qIviF
y9U0VWi3QCFaYqeupXP6fKsQHpiXVnZoUh/tpRVuLu31XUrOQellfz68iinWRfnm
aVdsJXDja8WzIwDwIZIQNQTDYDAj1y5+hMfVpJn1I1xE2qXRI11eCCJncEZfr5dQ
rInNBoG8uVP8myGUw5xSwW/W+Ckuxe9fXYoBEsMJxYrrgudo7Qcf0FmK0Gy2UtUO
OuRQ5AFm1k+zGvAsfL0QF+jRrQJgKIYgNuH2kSHvzzoTVJxNUxoUpeYsV/JGrAE/
7eiuwoFJemYD7R2e7p04dbITVbmYnKxKgw1UdBf7azGV0qAlH/6vcXNWhNupBHdL
9wRThQSrNdgi+3cqbiPwgLu23dL6KL9D6ml649e+0h5d2gp1P275IDH5F5ljNr76
t3WFnfeq3Td//CIo63ktSQL5wLQNLt3GGaa80W91f2qtsWqr9Iczx7d8+wxh9ozu
1PWANj75R/WxXEO0CobVIGdIHxvtWx/sfVf+2vs8wlXBDPvTCb5KNilPkEs6j044
DXxNaTPUhAG2MZMGeWdtjx2mzFJV0gf6iAmlEyGqLv2h83YKfMgMup0eIMpcwaY+
TxgHngQUWieuRPGVi2Dhp07rmcJaYuEN9wyNBns0la2WiHiZ2ddC6XTJLjXuOB4x
x+4vow/YzoVwZ+wMJeL3C6/xFO/3xIzK6wN1QLTn5SLO+VeFrSaVbgVq3ZB1jnPa
8xM+EA6C3fUIs7C21CcKeguAnjr6Uo5cNBB8zNHa8m6LG1wM2B9CF6r3hjtExbaa
jseJ1BHKE/HrkmGGqMXEws88XQ4e5vn3yhlCxUzuAze/inljaA5hTt6uSLplQ/UG
2pVadWu3nfjn9cAMjp46zMCfkKhbxurV/e20CCMF9l0v1ruSOjrOk5f0PiRIUPzQ
yKVxQ51iwkHc0jDsRpDRL0yKtP26V71ELbaiuXbEPTSYsrBQ5B+vNh4e1VWxqI4j
U+c38+s7MhA8vy84LycXVUMYDhq8TiXG14QxKFMTn1bNF9QJEorKtjSRisydsB7w
31Psm143DXS5zs2ges44gcruf2tfXCdoZby0BFX3RXzU9je2Om6NNeQA4qiKy0cu
BkvrBJdI0A/VA31ZLx+M37SUK7CSjZmyKsXa0U9zceQ6r674ReUz+wMzjH69FRXb
3BB2Mqc8hYv05Oe+MwC206wSu5BzKQUtqBzsVP+uc6iKCbxZFZStho8MnCJFdDR4
HOk3jpQuj4PfVzcD4uk1vgwCWF2Q2261xbmfJnRNwYOQdt0SPFcVkshmsPO+KpYp
1UQWXN2xqpZhrZk7R5mSH6gCYLsIQkm0HPppcK6BsPE4X5m/ftV5HEu0cYC+jZNs
xHEYjdVWkRTU6iQ9F9SYRAThXTmd5mdXrymkwTYtK0EFta/MAv9EHRFVxTDHomjV
HmJzh2Y5Gz2n/yZDUc/fjePY5DSQD3ec4F1NahfMtNjNBwbAf1Oh0d6bx9yr40Kb
8EoIxSJ+Hcl90k5Wl4y/4tA89PFHxmZoSqJ1RxajGi/krQ4vrjfX6FDDsQaWg5by
lduuexBGLHjIq4+RGUOP1r5L80PHlo3mNvYW4g1n4gLycR+rOYxVeFMd5dVV4NIl
uAxTKL91GKx1zhFUQYROaZyFOwxF+TCOVYUHjGR4PvXhiyEgMemB67MwIh27Q8LM
O0pqMfGp33YDIbenR6JakTUPLbDzSgkrakRgyhyMmeawnXj3qGdTa7iDLqS6sCb/
GCEwh7FB+qPwZwzyml7b2/AX6bVwUK9CcU3yNB1Xlb6z0jqxLbB4+3bepcas0U5U
zMeenY4b3KCpk4yaEKXD7Yj9vSnIYGTEnM3tvZOS/nXOLP6WyYpR0NoFZEhg9ecp
ts4/3wD6oQlzvyWsgXIFa0cDobbGDxQf8LQis85Dkxb8kTiZqfruR3PU0usyFI9j
o1g+sckfX+X7g8QRakt7c6KcV+37P6YTSEGqs9VLon/UjpDS2ogCckVexHa0XIny
3WQVHD/blorFIAz8JVcZ9vdzUSk0xiZ0IMPU8nXnxWA+/V8OdtUDx7qqWFof3ICc
IRUo5fYKAB/heyiP5JCm7lmU+4sswnJip9ZNdI0314RWXcb7tEzUgKxHk40GwdxK
XQCr6zFxE7GDKdqXwCXsAwnGX/Sl50vsJQM2G6eQIPfkKz10M0Ruif9lZKOjChC5
+0FJUYoalci7oULevnmXaVc4cCKWU0xWKldGnKGpdsyg1IJsx2Gi1XjLAiBPWe1d
WoGnIaDG8niLf6E2tPvuKQr0pM/D4qAHj1WxIAEU5FgRE+abnkG/yKPECL8NJMgc
edTi7slpCi9VrA3tAzR/qqY2uS1wkEy0XrZKCk256jKrnirlp0s+g10R7zqaCz9e
w/A1y4+R9QQ91b9On1pMepp0KXA4sqU0PxCtmUnBgDpkn2H7mcNj2sZXmyGMs4K3
uVG81onsvMvfonlpvhHSsmM61/3lca6PUBdz2acbksdGG9o5wS1OomrUv7BL5oWL
s4N90kjvwLfND77b32zpGgTreQn5wGAwOOE57dOg6SdOA33NG3eHK7laBn2NDmZC
OyvgOXd4Z1djJJNKsOvF385hAfH3E/ASNNaU/FpNAYAxZVv80QqiVGjdrxRtBhfy
Ic0Vyk5ADCNiPvRUaYSJP/vHTugklsFxI3ZTCrAbIZdyWoGvY0E9fUZ7obqSurNj
qfBsU/8Wxf8c0gL/EaV/SybsjC6mfKVwe/oFHIg3nwityX8I3labMRD6bQKmMo9O
Y/9tXGIzu2iaflKqlxFL+dnxiw0isrA308EqS+llGFExCFk7zpwHJptjbBpqr021
JjOsWCo3FuqBJHsAhu08icfEWlBCFDpMSgyZMyuE/qsG1vnmRzXbZp6FrPL7tfio
ohTpLHMY0wdUfZWJBBbvNUELoZLRfmALVqC/ZZVBprjeDOCwWjqEY9JzYFDwuWCo
0PAE5HUhvGEuF8opuSyzdr6tfi/eXE/qoNe4Fs6PWqoc4bqNvsfOIHs+pn91NGoW
q2NujsS19jc8mZpGJbkX9qAqAGoyZMstuJXLTyAouYDMlTjg9vOGrnHiC+AT8JIv
zEx+B0LcMapUb/ZRFkTjJlTwrmXWzBBI7SUxndoNkfkzlsXCARq173igrCpvO3gv
2sXaFnbJkMOu3aiZbqAkmyi3kk1jRjyyW8KT309KZ53WFO9pKt0NkaSMOK5t0lUJ
JCWpKbAbvF4zYnfZWt/4whFoKDnEfxStxioKuPwejQ5fA+qilcvMOLlv7NMSeDpS
kpaU2jWahtpNpbm6HenheOpyZnEop1cfwtLcCq0fiMfGYP072+3x/DxcvXa/JbJY
wmfcVbYbXHzLowJw6xuNVXaIJysoyRsMmm6PbAVKu0P7ysqbQfiHel4zHeED6P8C
Eh9UsFeHlDX40D9e2xIEUb0lKoRkBaRXLUwzsj6ZOWLr3bwsr/hCgPDGBHK0BjjL
fQC/AbWj9bJHfoY22jhAYsmlZL3WYZuOtdHDkA6k2XMLgyieLo+8/mZ5vF7XJT98
zGYaexZXSbNPGXpeyns0/vI+DY0ykRSC9j1GPSjlpxexgbp9VeGwhZADS6iLr3aS
jbuTie8s4P5zgGi04ENhCjmUTwaYBb84RBLZJoBbAbdd9ka+9dDZDQ/zT8LLfAhl
Ifc7P9On/lNhVdcAAx1BQMxg/EqvFyR32cY8rWT429pin7UaAUU/m6qgVmuJpnJ+
KWjATSKGQtDjBBMRR/LfOZccUNF/EY/wipFOq64nfUut2A13nCOJrckiP0/ysaAZ
eYiST1bsGLBoI2JaZIg5jJErGykwrB/mKKxCeyKjV0A++pt2NPnqCsR9jOQQy5bN
hGykPtyEJEwOiSoblLA8KtH5aUqQF6MgU8O8+xTlMMIIf8jSNNgdxU4rU8uFwLkD
m2lSQ16Z8ffEF8z7j0HXpT/ndlIkZAs04HHXiYkglawEbVRGrBq+zDQkqcpZZ63d
FObX8z4LTDpt9SNjRKeDtngc3s2rpDYKhQ9ZidTWO6w68aZ8T295op5gaSxLhyZL
PRMGHVNwJ+tshbC2BS5JBENUBFR0hE4m2/eCGARHUoqxajh8InRVFO35gTrhxTZX
yzTmK3YeL9Y5I36IYzcoSAVcjxsnjlsNR/I8TIt6OW5Qyjn9Eyen2mZ2lpbEYycr
fznlhchTZilIpo5cSWkXB1klnhpEq+l5qPeO9BL8lJ3vp+twnC2+CarBj8XrbXWO
glkrcQy3/czs27uRVEcnCpj+EoDHKo2/29K+milZvtqXg105qOL27DEgarYrCpeg
eeMriveA8OF4X4wSgInM9XZazGyagysT3u8VCMd5DDCgh2+pSR0Hbeeou2TinbgQ
4lC2qAkbLzUYfuVpn3Wnm1ykiyfYG/UUM9XqW22spHCt4SoYRSi99Cb37QDb3vzX
5kgaTBYDTYhEHF7TtnBx7FIargUnF/lhvdgAv8CQFPrqz44lUSG1i5FJ5/xruXmG
bL6sB7dcC/DAPObzwmUU9pfDRpgwcrWoQ06jFsVulqSiDl9NWsn4uUhy36EuyPnR
U/sOTbYuULXOq/INaNpfud4AjD3/w7hAZER9+5JbE3nRFLh9kK6O+E2mawTnQZRH
dqanCvQ2S0lEeNoay6pXgVCaxstjQUyTkCpNx8OVsM80g7AOHuEE2tBSaCqDC7pT
AP0YCbSXtBEuYnEoNKsnIwUjwJev12LjxSM/oZUzW4GllRse6V5VvUHKs2yeoAfV
q0IlOBePV7PtiF7UggU1ge2hVvltt3pPHwqO39ts5y6HH/huVcnTLarmmCWPT9K0
8F1qcKy3B3qZi6uOj/WAcMBMKZp5/z0WWx0U7jAjSjxyZd9TiNZUZfDUwjyPWBT7
xaJe5JYGpGYUjl47PyHbmmqqJH3s28hcGXCXVy/J4OOvkSQj7f2f0HQmUgT1MYcB
XvJYw1ONOfP1XGFlL0PHAWF2+baHP7Se9h9KtWiV38fQPCRhrr1BeXU13EeaSIN+
bzneHdoduLsmYO564VLaCJudDhJMGVhWaTzw5RB0r5kqbB70piJn03zWFGYiZZ9Z
F5NN8suz567RVyiClgLlRcHje5mRi3lkJ7bbcu1JQXh7PvWmm0D6MQqsog3M0xMT
wIf+lyeKELPH5KIwPuQ5QS7VllZMC2hoIK9QymOvRQY5njadV1aybGi+RW43dKJa
qSY6cz9QIh/tPBC2QfKfGGDjrHzewxdMuu96owrCdHjXLKzI/uNJR90qnKBZGi3a
DrNDIwOiGJxKWHIeNmZn93FhoxIUH1xiuV5GiIuyHoMdNeBgoF8x/qUxHn10C+6k
hKm3+F8DiSUV7f6dEhdkuUUj0IY1TY8fweo3jM0sy6QkOWsIiArmqWIM/B/ohoBA
B6//TunvTpQertQfYRdfwkXPDP56nwrQ/xgeUGr5k6EaBysdx2/WOcMAHJ61w5rY
qPKVy5vNKABXUZqmWEF3gIUv9jWPGJcsbKFc6Q6Kl+66a8NDrXVB7fGlXv/LIDF5
Hl4xg7wAGt/Q3QfVSLXO0/hcXLMcHkMgHHH7QbYsrCCcOAv4FknofiJK40/Qp0f+
J5y1n1llEMfpSnDGNbamJityfhpcQ3qoOb8mJ9jzWEgGc10JYaRL+ETkAnddy1AF
EYQMN9usafc46a/UKG/P4WEGiEvavzWwZ+HsVVlpfl7quB8JktlFHOMC2tb7yZI8
pI1U+cIk/SIj8PMQwasTNrAJ/9EZXBfDX/d3ZBNmWhnJbLjeu9SWjkcYfGT3Sm2p
WXuFfnfsBoZrhqnAiiWVAzwwAtwPqfCDL6H1oTqtPoszygXtLuv65qN/R5ZCTrSq
8qi8L3Jx8aVtvQyo7t9PH6pfNI62k8t+J7OKj5hL8m8kAMWd1Tqv9LRAZ2ry3ikT
8Ds/kUH574/CnVDY+dfD7q1PDhZ3d43rMfFBTsXDkYzT6D5/tRtm1eeQ2xvC9wJB
g4ceTA/20c3Rthw76UJA0lCzbAL+HUjz7zKWwhtn00FuuC3fvLRO9WrCHFQIhLdC
nDeFv/H628uSM+HxTyiBGKBmTEpuESGFqQnFG5xvP2qrKK3WryBSidUZM2UDtpaO
9J2bmZ5yIBe+TXGoyiE3New7JIsRR+AMa+Gf7KtW0tmOFBsEgdt04JvP3k1yb2NW
8ruGajGhofH1LjNjia4etIm9WNsyCUZxq729szKlC5JmRHr49TC//BcYPX5Ax48q
l6vBnkvlW5VSfpaAUBEwHlpCbBoW7IwbHcYl0uCQQR/w1/9mRt7er0elXtnq8pa3
qKkZ+wRBQenxBoPAyfjBHVU02L6IhQCkBVKbpPRqeUw4I7TPMupzmyfCpKOmOhs5
hy85Rfp9DsnxHUxi+Jkvhhx2T9VvyYvaZk+5prllKxQoanZ9XDyLc8vC5jo5Krm7
fQVw8FxWTOBkRhMtriGQ96xYfTEYwiWxxtC5Yk4cJuoQ2XCan9zWoyP2E4nnZTJK
PqVJM8BxSfv31+wdagl7rPRK7XAlv1i50PW5wTbHBTYJcI7jhIHJHHtuEGCFOeVK
o0/qlnPzyUsLvhu6DAK3aZjOKSrVtGZZSV4iGeRsaOtkIA+AkA1Z4kjAQO0P02hU
smhF+Ni+wEEQV09Sg3Jdk2LBkvfDvdM7eGvATkNM9aAqNm+MoBxdNBa4gFT4oTjo
9o4+y1m1cALSSwPVtKilmNir+M4luNiAIlsMPdZcZyyfkS3F1SurN8HQCPf3jaVi
LHbS9B8sPrqoqg6rzFTfgh/dIja4M+Eyj32mg7CcIA++QDwsFPIovN3+pfZl8O88
wbkiBY93XlzA1eIEE7HDWRFuBRNBTyZ2K7OY3VydZm/IXFIBVuo9VM2r3AFHg+Qq
VsQxR1bIhj68BhwcrYok9TnNrZW0elnwP1XB36DYXnH0PLIqgTdLrsfkJ2r6zUiI
Bgp1pWu4ajxYwk2d/qtUoCcnYN4eiGYilFaikb9hTQAFogwmPUaCyPz6W11rT/Fs
EqXmICq2BWgZmR3GKvGo56gs3pzdNxDC5oo4t/CKWP+4/wbD5BEPkKTDqBsibAIK
q2HuHgVl+/LDiGKXLAA/Q7JwUB01LLLkzSARK16IRyD/VllAzddI8rOSfz239tI4
+nPt1izNu1XhdreW9vy3GPywCEN2WQ8ZprI8HzDhUOtVNcHRMBCult/pblwv/HB0
2cX55tVJxI+6W4JJmdEQnbov/bUcYE74/exIxg5jaKkv/Q2pmcaEms26eTOijwFp
qfkFim2w2jSKyLIP8l0R0Qmlybrndz+/7ahQIyv4Df+gQvL45wvnR6NmwdTqQHzh
Omm7XEjWiXIj7RYJGgIzdhZTcI2BjnEKIMZRdrkMw/7HwCfCjXKxVJsDAh2DWCqr
gCfJ12TJIZCiP6l9yuYgjZKmUkmeG1n0M4GFeR5EeFHPRMlbh+NeDc/fInCUN13u
mtAIo9h8N2+xSD6qwl6kstBrj6st5Et0IGVAUg/8wkUsOs4LX9p2KLJlappCoZXc
E1QkFxwk/1drdR9HD6jGzvdf9jyYhSroOr2vw74fHBmTQnP15O2cy4gYyk4/Ly4r
4rfLqrP5S9igVsA9AXqCHtstdtf4ywvQPrn//WuRe0eVJlIAAfFaQp38KnbK8OzD
UU8u1sY9TsXiv2dSNB2gUGcuP4aicQvyOGGNC/AMP0icdz4EtV1yJJzATOYI8Gi8
1QlpFKHha5n3NMVTMTSaPHtGBa+XX9TAN1VfnFEbcnX/xu++0iuPVCg2cVlqPBya
WKNCAzwLY/LBfTT7I4uhuJN4eReCaG+3MmKot2RJzZSgA0NrJN1dcpf8ccEhZ9XM
bHyK4BFGr5jN92NIu1KpM8IeU1PofVimLpBDwUriBTA4BKMf8xLTUVZ2JV/hDGnh
MLxct+9d69v9D2UuhZV+DGD0nupiYOclYjzPf0VFm1aFe1pATCySQQe7wGg1eeJA
DqUMVhHtRlLJCfA5rNsXjtep1VVC8Get4NZL4icS+CKBwff++Jca4jlLRX98d8uk
ZqLhLKSHnAqxDCe+ISuSdD7wWLbzGaPk4XF1wMjm7PoRCvOnGFfSQ3TXXd3Bc/Qm
STBrR32s+vZ+14gKaw7H4DqX+IFtzyfMy53sRxsxZOHP65tF8JbR1l3Aw6CJN95Q
ENe4E66GkkTzkp04VjAIKg3lEJaglZvcIzoaaP90OvzfitFXF6vy0cIxbIIaL+SJ
y7h1yx2Vz23mFuTXH9E13mQJEQC+ZiS4GAyGoAa849JKyUdnA5wUS/IpapFAYYaV
aHBT3U/J8q/vI1VFpoykyyindLQHDB39LAm8QF7h9MJZtpeJw5y3NLErhbHDeN5Z
WulSM15pQ4d8y6t9joR7HQcaJcfvTCMu7PZcqS8AlYG61CH3FDaCaO251zwk1co8
dnfL9evqSdOsaVzzp6HlhdqI50kTBVOmabH24oH2qS62jOR5JIgGud8BBR/uoisP
Q8CezkQFVICN+HalEN0rmZne/iGxoc/g/gv88wbSC8IOuiMIpACpB4gxGvHeXqDf
HarsvigJVGYLBKKt9BBckJWxUHfjda74UUoky+cmD0jO8fwQ+aND4leN9ThTbOqm
EO0nrkd8Y6WinAzOVvMS5AUdOmxt2GzGjqPeekXZlT/MhJHX9rhdMEo8VB+SkXAt
IQrpr0/W2rdjW649khiN/p0/QyvwSxP5UITxEcNsD5vXgdBvF7vgJhEmu7g86Nw/
7ghZlWHyXaUDsUiqKZRMJ5e5CMSv+fogpoP1kKyZYi03RKktHpF84iHVLJj6dGtM
gWSNC1t9oMNO9LawatGCo/lF+S2UJqkIJEuNlcYj84GpQ1inEfzF+B6xDkJELuiG
xf7tYeO4ue1+PTlVSCNVemxesYuDPa/75bYC3HJmx7CtMjFDvaP2xIhNp9v99xZu
sO3jG6itT3J4ED63o97u6BeRpp//rve370tPcBtWh20=
`pragma protect end_protected

`endif // `ifndef _VSL_SBE_TYPED_SV_


