//----------------------------------------------------------------------
/**
 * @file vpr_intf_hndlr.sv
 * @brief Defines VPR Interface Handler abstract class.
 */
/*
 * Copyright (C) 2009-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VPR_INTF_HNDLR_SV_
`define _VPR_INTF_HNDLR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
DzmoCygPEYXhMVh+Uc/ZxNnpvos3XOLp5NXEc9N1zLV1n3H8kERKwZoBO6ub6zRd
Qg5Yb9F2CKsdWXFC/NUZnbVPmH9+q+qBs32GgaZPrTEmpqmwIOV3YuAcQLpnVWns
OGSvTeOXM5SxAkHOfBaKyit3tAxkcT1txJOLVPdx7dm162qdQPBrqaODc/MO+M02
37vgGKSSzsAiWCmtC6NNEsS7LmPvYYyIqc1k1aeRcoJimxSBhPC14DI6jS3udXwi
779jWZpNyUhBc+cq5ePcpPGgH2yRIsWWtsG4M8aCIWnSURN9aHPwtwjHLV7SVTU/
6KT3kzIG16LTq4pU2B7Gkg==
`pragma protect data_block
4qZRBZ9ygEvGch/xUmaC7D8zV4axJp/epM0EBdI6/OP1X91sUsRqsxpV4fuDZTRn
oun8UVcmett26hXvUHSQPf2V6E5Zp2NnNONWrn9R7W8nsLlhGMOuuhMOFaTkhRwh
g+VlGv9Pzqxykzm7jxlZNsiCaf+LQ2Slyu0cXxyoFAFY9uR6qOMuWyE2nqRcJzgx
HD/KPNlBSNZyLT1bTfBWitDJpYU+oHrjff1SQj4pl/OgozJJCTE/O+6Pfrc7W8R8
aV4wFRtrhw1xQHJa1PdcwZm4dtIi52qhLWYyoKtpegj9zhHJrrhz8aJ+ktqgFJvS
rG1cheCHx/udJ5PlO2Yn1XPP4l9QiHKiicvIKDp3ANhFuwqc14tGtv0XtPJFsylC
PU+ZQuNnQA0kWhG5o9TZ4khIaOqEbbKypy0V7HL38OcpyWCSjvpoNC/B32QuuhyM
RY+TmPhGS8nDMPVKiJ3OR2cV94woddcVLYOyJ39AJ7ngHYY5NbC9sSG+QV7dbZH3
yyWiOFKex7ycPcZ8cbm13W/Kg/WgYPlOPigPiXxtcDhpv03C36596Ot8nXKaJPPx
hVGwRCpIo+mlUfnJWdrRRn9Lfcp/9egKaldn7PlfjY87XnOYjQjQ4fwLReE39T7H
2ZZgLWxbJezzg08JN6Oez/GoomQvZH6p3AlGIO7cgMYQ5GD6g3oa2P7+WRDoa8yB
/156A39wwcLlWbJemF368MHpnNNMq2/jtq75RMPENpfOYn+BTtpMNdluRmyNZ6we
4LWaNXFUyIsabJYbrOgr7GzR4M/MUCx4rJ/YrdMmzPPzvhQivIcYOzW67klb1nWR
A1BBo6BxGZPZR68swUFuQmr9OewYn+JYqEs+46RfUjX9W2KVTnUJETFrDmAYlxNk
8KURa+h50ujSClVXXRZAgwY9xgWm3amuhRbj82bi3lxwlBxO4krAgzuvHGu2Jg+B
LcNkST7It6XVwE1lHygp9oHX32/nqJMzY//E9tIvFtV+prSlX5EAQ2cfWZ/P58hG
w5cpKUbK7Rky0tp1WjcVAEqGlrdg2an766ZHeaCbVhQPOlOkCTcurooBax2BDayP
fzeoYpzJRP+imhxqad1o4GrmSCQcu66W/JbhAw8wzDppofjfjoen3epr7OY2U4NI
DpQ/C22TXhJxEfUuz9PYW60SmR9BJwi+SQjVMTrcSHNs5OywncWSWs3sVGFLgphG
/ZY1NWA7/8m/OZurqQ3ygDDxUn0KW2WygQxzQRMfbFOBWZl9ua4BNmhNXW1O2AWu
7KYXWIUea06omlCwk5mfc6it9IGGNW+ljexlKVfAGkSJvAfIkHcAbNTLs5SWUxSt
JdOOiytBAg15jBUh593MhlVisrfTJXBTLlad2pI5UCDuIutwyU68h+bfOH4Zsdcq
6KBxI40H1VyOzntO1dgSDD+dEWodJlzXWBRMcEK+32WosrLLadj6QHnlJu316MjT
xuQnWYrHy+QkAIb9MpWYkdoaCqp0UvSswqlCAGyOEfUg3debDP71mwLX4e53qHwd
r+pPcLb+WdsE1STyEnxd1eR2fJglUxD0qfaf6ttEPKUcm9dfQFWhBFaUNgitr5ku
JwdjTKRazZIcclSIl/YD3Rqo2uufkYV1ZW8k2hgYsNb26lprfhxZzNeCBF6u2jHv
a5VhUNsH52gOYwq2XtTJDzkn7VJxJviS47g/yaYe3C9xSumEjgLvaXkdsCz/q043
O3X0rMIUHJvzy7NTMlBszetsQKjWagKDQEsFEAO+mRdAZdxG0ydp8MbE0EQ5m6KV
SzfzlpZ9eWkbI8wx4GFza+egjAfaLkbLWfw4f0qVw+2AKpNNd5XQgBAGUBc44zO5
OMMxX8+ScWiox08SNZwL6lHX+WKFLSrQ2R2OSNQ55mYxJG4NNvVD6u46VBo3t3zm
6KTmdQoo8uhDACEOGgx1gRBLkZIUtespQn2s7zZFo9DAjQ/HEdnL6rMj0oDxspYJ
TskdopUwyVrA6U6LBydCqErwHUo8XrVyGWjUDl964GuytzVCln40ES0yXY2POaSV
f4DwRAiXAFQZJ+vPs2NyM6Mic/YU8ULO8zshao2nr1WobrPYXHjSIiY4zvgZ5eTB
nKmfZRkopNCHL0QM97wRZ14vQOXBO+FAkRNE1dgz9aSt7tpSCzymC+MBMuUq8r/F
y39ffRLpE3gsGKUZWyIuCGKaA4j5D5x5CqDLi/ENNsgQ0oUONBu+G58fmpGCBK4B
lzlDoDlcthuHsVKNGl4IivbifyMudllkDZBR/ZimwwG2mI2Wy5DNoVYhCHn4/Et7
CKQ2DgeCBYCsMtOzgR0dUdMAq43l9Yg6U9/4aYxmQegMSvSwKXnP15fnhy2soflm
PYqJPFgzbXYHyIZk/kbSET13IY6v1H00Kmft1MakDa59ga1606lcGPWB/w2GeV+9
9/7n6DQ0ZbSqMi4beBnSoRmmiUaazqxPhE0rVCx6c3G0NYsG+dp8GRGFllMOMBWQ
To6I6N+rdbS6wfoGZIFsXv3flOtkYxjBPCI7MBfAAfvgY1Ol8xrA1djvaVx3YPIz
obF9D6W+Na7MG5cvOh7DPDPW0BdvaNqJDYE3MoEAiNitAk8dwlm6e8aoRLUNUboR
grCmFkoefcLWNGAfyq057objjlUMbDU0A6WPVJQv7D4WbKfCeX1yHkA5djKRkmJO
6GuUYUAWr3Usn2XoYcXiMDz9ETL8BWR3E73W6Oud60cq/XLjAcuLcCLPNp4B4M16
j3TFIXTXLveTGI3yWir37CooaecYSBOB5RuoY3I0GU2ZvxLFEGYzM9klBdtvVrba
2Fi7hMBao6tbwJFMkBGllSCeIA5vzoAWGrA2ZVthzID1MJA/6qxdzV+xjCIWYdGy
/Zu353qEbttsOs/ubNM/trvOZpteyjxTolhAN9YgczW7wBkZ4fvmGA5k7qOycU5k
2wnGQNhNa6O25H6mjcrKV+ocL6Z0yYT8Z16oFDJbL6VXofW2GevgNBTbIu2na2sc
THt88htxDvs2YJ2zbGolI4K4NKKx3XQS10bevttDUAw5cEHX54Xy5Q8pEtqDoNFH
Zoe8VNBM0/YAPIxaS+L/iwDloD+Qkfne4BLBhuCkhgTSArOPAtLKS66eUHtaWLra
xew/SB0kHc+lCL8MRAS0sb9kkuzkf4l6l7qR/Du+RJnxXJDawiOuNL0gI/FqZ7VL
G/S2IZQAYrUdArANr+jyDd94tTJwHo3WCY65Q57R8KpkoV4If+XCQR8AzoPV+h6G
kFMyzrgFJw/mkeFRqADQoUChf2PAQf2xP/FwXwB2uRfsKH926xbKXiqbA0NMYFjz
Otl4zF8N8E6sU5AbgOh+r+Zn+jx57dcBfR31orez+7mpiGvxf2smBOztHfKKsqol
VXhbfzdiqiddxwJrAQLq58b32BxRiwscvJ7eDDXYWOY2H68maasnOQX6sgiY7GFH
QHqUVNEiK7JVKxNMF73GyFOtmIuHc8lifDx14eDkZfhEaBFlJoOnFwXHKd1pA1dg
xhyMFO/EY2aQ6H74s7Xf65BK7XEcXm2ehlzXhJBMb5qykdJWqOEGedMYVXYEZdA9
SSGdxOci7TstFPctrH7S7SBCDLvog7MtKBtN5J9S0NkoGq8gOh7BxRg4MViK8yMu
ZXhWZlaji5/BSBInmEkYQDgov1ImX+UFbBmiM7aOa2A8jevZvAea3vrB5oaNqktk
VLXfkq1whE/gxmUgplPgcbS0Y+Zp31WK9WOExxCXmwHtdiuNH93dEpu7dclCXakL
HJRytcAYjCRqZFS/m6IP2ag+oynoxxMdRzQB+9JTOZIHAQxbAtrawwCBrvCpl0Ya
V6JYSf/Tu8jNPaXtpH0/HIswFkT+HzrqYQ7zHG6mAAS+DbVxD26srUk1vRgcSn44
kj5jBWw+6BNiwn/mt4OJ5CrQJcSNuTqbHZo9uSO52fvaWhe2EIgculLuT19eEDw/
VOR9Ti/J8mt17zcWhwADiXUv8uLIU0iK9oNEg0wklr5ZMfY5mCTzVOTLkP2Fo9S1
f4YyJvZPh4Vhy+5i74dQYe9wTBbMjgeA0PtrdUR73edi/hRvbVs/set/n3+NShUp
CTLEsAcUePXqyuZ2hM6y1XXEgVRMDXwlmvvuJjQZJoe2edSjrpO2AgBx+nrEkr5c
YAZp+c1Hk4Jrt0qofJI6klYe3dwDDko9EldBynAf02GyYKnK7vOoHnCLLOnuxSPr
srN81H5LtbjUB5CLY//9Hf1rBfUfhao4Xbd+3u+AqBFpTQDShAw8xUfTFCrS3WbW
Wiy47fih51B3PbEY4CWl82MPKmzfV2uxLsUbbul5g0Ga4rqdVtsyVdVb0XJ5+ZjC
uAFeq34j/25A2ggy8B+bAFN19LMOmrPNovh5LuImBZAscVenqSeVR02sSncEaulg
v1HTwnPBoH79WpretW5hH5oC+JuBlppXkwFB39FHy6tV1eIn9mW4pT9W2aq3ZLyQ
s/jqFwykdH4gWMpvk8Cs3bbZCvT+hIIVoAYPIBMcPRPowsi7ZTvx0aVXhqiz+ECu
9yCPL2CILxKlMBMPFAARXYlyebhZRqQBM6OaESgJze2HBO6/X4AtMhP6I9Sjr9rn
vZRpwGsEtkaiJ1S1EsoTnDRBHJupWQJKDKFQiJB/gLgWbY6YWesBZEgt6Sl795oH
3b+9W1sXrRagglx8IDeUt7l9RjLwOYeyocCRqFYjYELQdd4mz9xS6QvwVS+ZiWFv
s4r3DNYJBdad1rA7oahfy1gpFFWd036CDIu2U99x2ZwNtSujyhlHYdiQQoWGHvD1
VhkhMidjm8u4ligwkUwZE+8qotskE9QasvBI2LW9xu9Ay+cxcG/lkt1p5LwpWJHv
aq5cPB/L7zRUk1vT8pQ66XIecdF4h5JL/T0RWl74oRvWm0srsp/0nOg1Z2nb0EmH
wAoh4ryAEZ7mFxGaRdZTBNiaTdc+7JrB0JrtwzvkjD5OCWY4hLOW4oulxaf63bRT
qdL8WTWQoLY5WHnH2wD1yHG7hnhWusXy0zMd5P/asyTVA2XfYtJdmjHuiSKIF9Uz
O5+a+pXjG0Xap/HTsFKjlcPD7iCjD9SGGspWIurK1zp8gUDPY+uRPBHE0mD2zKaD
mLN8VSrlGteJYpSRFq5PILdR9Z+goDUf8MzVAQt88cj2vk6MtxMjdC4cZdNljnV2
80E7mugiJOGDYglgbeSXxhIvZPEAQRJn+wK97Ai2bjaXzcwSPrkr/VUerw+DktAr
w4KIkhYrL0tOukAFVHLlKLgcfmLU/mHhn+LHMeSrqnxRebFxKvCV8G/JOYaEkvtz
TDsfJwXnF3AalUR9gFB3Qnl2TfdLflZz5H4ZPqMprZ+h5SGwbTTf8FeDR02TQoOo
lbUD7uqDE+ENzi1KOLJZZ0ZuiDdEXlArZo76QY2kiTpwhADPcHFf4wJYf8ISq5+r
Fdt3pdKgFflvPZ4N3+A18H9xtYqs+vSlD4HtUywNuNbLl9KULMElWLBhdBRCH91X
osyoxJiV8xlG5nufLp/jYpynVqo7Ofbzht7YspuscE1+ElOe/x4fGtkRAvwgjCYI
OxQ0NwiemZgYctooYeSGrII4UmaQzEsxZ10eDYCAPdEf0LVg0RXjAtjHAVaENC9P
M4cQK103M7Cskid6AWIH71t4Ia9hjPwVAgVHhD9cX9OPHMYZ4fj0lMwUQF9XsQv2
zUNbRcEAg8tZC3Gb15Cyaf3zwoxWtkMwZse47bRApxUAUgDsfPLeWG01Gj2+mZ5K
emX4c4MhDBiNhgbEqVFy2ddF0tVVtV8Od0K/2SMzKLyZqBIMGpHAnGqpkr0KPDRz
lkIJQ4s0386K4VfkNGezLF7JpYWXV5TVLByIQRoNXh+NAlzMXdBwbl+/8ZNLyv2M
Rje2QMhfVzSfA3FHWmmpvfQ+6JIzUvgPv36E0kcIScw7tKWx+N+YSjABwTMDFD/P
nitcb+ykgPWFfvrBH6r0kXo0476Bv/3DARLblsh5StAmDiGrkatkqjTzEOoytm5f
8Sg5O5Z7QRyID7Uezcl0ew1CBO83ExWPMFu4Y4d8d8HI09cMsreVF4esN/RKpv7R
K/cOkqVYioyNHBA6YhdkRb7au4vfjcwhNIwLTBpa4oET68WLiuo4ql41R2WrqtFL
gLMDuYuLkSAunFNttTA6zBfUVJUX9jAgNOaXytdlBmXgj5L6n8r7S5VMFS4gjImj
J82fvjhDTeEK/NtN+TxMqzfnVJTyjkQr1JOnGIullL6ZYd2zvoWymuEcHBW++cYM
cVJQGixodwTmnJD8elEifP+llATH+2lWzVuNuUDdWDg3fzl7j9kDPqbeeMxZULmC
G/B0+YqgqMf4QQe9bZcaEvQKDBGg6HfWuehAX1JUZNMKvz3r8ccOIa4O9iCfx3mw
QyLWOK918r7CHaTS26G472WArP3Ow2lttuGunKj+4xgoUZxH3JRYOWMGrylNmh+7
m4xWOCrmcEziuxi0sy1OJUcfYT2WvnBm6qCLA+fXKLHGvht0Cp2mAfPCB20l9JX0
Q6RgpTZ1DjRJne6X6vrJyhxGUL7cg3NOtHKDcXCvG1j6t3GN+RuDOtvy9+JOuOof
ejiA0pF/UX82PjotySxSwV9lJ5PSntpyZ3nawa/M3BMn5ojwztmTOTH4b+7JRQPz
+/ijkD78FW6pdQ/oh1+xfu6/28mW4UrlrKcXrHq7ZuVtDMIjr+L06HfrXs4PqOjP
OGDByjCHsOmDUm5yztzLoSf1fQjyN1LmC2Zz99w6GYql4CyrV3AWy++XX5DmvF2t
eRcmkRCUMAOaf9TiPSKRDoFEVGhpPc0u8w0hzqMoiMN5qmWWcgD3Se+hAsbl9vTw
jqtracvFxndUfiEUtf88BczHfUHIHWgEmRUr+jWiR8M3qks9JyrvZhcZw5yLggwI
4w2yoQihnj5hlZsQt6zV/leLGmfonLmjKSLxRK8+bv2l6J97TpL+KJXBEcOJEsLn
DLCQkOECb3dxxJTzNyDOfE+K4hWkd1UGaZDwswnqwaq/9zo6TXgeu2FnqPxx/t3A
qYEOVNwRJ8r02gZFC9gecntPUQ/qHrK/y8GssXHWyaqEvzxhBkA5knvF+ygKfphS
JFUKDw/WGnvjvtaUu8kfL66ui/NkQTvgAP86KLjc7YGpcRAKfXaBshYPxf1VRluZ
zMFqIJOLv0vxYw3hGvbPNziFRNN9K4DEisQeR/1F71P4bojGJwqvsgkx03O8G7d6
292WwELnlMMpPe2v/ARsZZWC8MV2jjYGGEcuOfkAW+K2ddilztaNlj/O7cyXi5et
4Jo72CEmHoOZXSWbX2U3UNpxwAe17RySclAdmzKY1wkenYqVsJZygYArD/WPPZKT
iM/d146OP4IxQbq7UN0Ckcf48Xmn9A29JZ2PJz5YH4wXhZ3PqA+HKMNfwL2hK+1F
wuvEK4u95NqhPPFbFCT8guCeiUj2wtUSKAL0ON5ckXto6iUI08qld9fRuLs+A2OA
9rKkrnTDF8cB71P1Bnd8kyTp6rEyfRv0vHutvpAJmT8TdOIdzc2eVfQlA673GgRO
1jAuyNf4QCPfuvhu2BpOxdBeehgEWGFoP6C22LzojpJnLyNou+RW66TaErYaCZmq
IZXqU4HM77ZlsI5ea2Zhj6bpLpMPSnf3bhndZQXKCLbGcf7X/eLYTvxasrLZBO/0
pGaI2tplI0IueF2YNEJTI1tL3JKbhtMdasiIEzCSB+YfLNeNIgSqauWtYd12RDJ3
AD0Y6q7yQZ5R99xtnDbGec8NYsKtdE/aVHhk2fYe0OZ2LX9o8BpVORRMo2fBf7id
PaDZqZqTe0+S7JxXzglLmkvKdwvLaZLcpVfeWlj2F/BqH0Xlyit0aEUENW3NgkzQ
6BiYQKlr80SsmaWhTBdWwz9YeKCigxtY51QR2t4tsM+ls4o+gw3XiQHcFr48NKmV
QbfOEdcoIiXhYfY9J0/XIuSC+XYSmFMZshdzdY0fOYRVIjwxotvvhNkHLJDjOoiP
jMmNfXX5MbLnLPK/HgAafC7Ep+4dfMizCnlYt+f6y5YarVt4fsDggxmayZncv8oT
/Cn59H4LH4o4yc61UiYYiPpTJkepMr0MXnax4hvKvUCrp2KCnGEoeIECZ0D3LOj0
+/EaW2DP1+Fa/7HDWbAOCAB8GewWFb4RNmHvooJP3sDbA4fWXKcQiStvWNb+4fL2
pShCux6CcFU+GmrtHCMAj4Fub1YHeRVpEpUWU8VEX7FrpXIDZf2V+zi6gnoCcfjq
KfZfCDE09TYXND1fZUDrWSSV0x8cvKZPRQ+qDwGCU45ib4t5IAGCR+/xqZn0qkkk
pcummDlHejCGhTFTziRgyR1LyGIv3u43dSjt+NxFkiHO+Nq8FNz5HTYbUQVEkBwk
N4x3EwhME3cgcsvxZpd88ZGla+D5a2IT8DPVHFyUQv7m2YUkiuSFtzP/6saK1oUx
9gvQ5VqH30hFPDk36gLkmOItCSMgd+fEnHvRuR/kcsiH5PtUdA10R+/ftvynyqOW
vxxAT52ivjufs4h7DzR2ZB6pGfF+LkJJhZDFrCfPuDwxDCBB0+KEd/k5E+mncNFZ
GR4tf/KZph+UKv+KJZTw1w==
`pragma protect end_protected

`endif // `ifndef _VPR_INTF_HNDLR_SV_


