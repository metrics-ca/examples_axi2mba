//----------------------------------------------------------------------
/**
 * @file vsl_addr_elect.sv
 * @brief Defines VSL address range election class.
 *
 * This file contains the following VSL address range election related classes.
 * - VSL address range election class
 */
/*
 * Copyright (C) 2007-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_ADDR_ELECT_SV_
`define _VSL_ADDR_ELECT_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
nBtHf/UETXh0eWhXP7L1LTTnnxJtY8b0RVsKr7WVlMMdO1jz3++0pMlmP/lY2IXl
e8fkrUypRaC13Y0jlLOxkVOFAj/LvRpZSgx8sUg/8Td1VEU0SCE7UFurShqfHk24
S7fgIh/OkClDJ/YC7Uwyj0fWXpyS5LuS3O5xxySxnY+ETYzkr86JugezLW13MKwu
grsj+pjp9bGcNAAuJbPAAjn2whxqECL48x6pCMXo9ikCQa6jKl0lICyXlrqOD9xI
BSbIlqsZpyX/mLT7I7tDK7FibqQ6T2S1dDUkq3MEiCPXdxbomaqe36pF76nFKgEC
dQrc1Ep1WyhFoq2K+jv/dg==
`pragma protect data_block
9H7cAgOUrQh8B3VBNQ4iqWw2FtvD0/cudi1SkKbBQllZ556y4wiEHSnlH4LN34OY
EMhmXhMi5wNlCZc9B2gsfN4i0E2pmHENCah/RmZrbse4JC+8OTSPEXG6tGuSAF4M
Po/FRDyQIslV5Tp/Uy7BT8cbCL5NOKGmpccmmIctT92+Jb7lX/3IbEaBfBi71fps
gINQ5a9oT2D99Uw4/wVkgU2bABPxX/7S3GdRXFgbXLkJ170tA0jPTDxG/kZz/4eT
aQJ/bXs9L/tXtTAtQHBHixqmRSw3CMegOntywWkvCWhleawURElkp2eeakHufNvS
I9gGZpFQGXI4jF9P0kGhgYiJrBSLaqng2dX56mbhPObDpq3qnkARhzZJ7HoNCMvb
cn4C3JN38PK63326CLAM36jUM5lYnHvHFLGi4aSGIzENmTTpCkmR2KN/85PMIpSc
TSekQ/Dg/SFbLnk01ZisKiTVDT2uGOB+hgjbI0cHRzpL+dQMgw2kOnmn0efUUdMX
3/rNJm4TxgkNZXfWTOIy7z1tSMbj7vicQOdn2AgFQ3g7PDXQVhDoAcdiiHnNdao0
nl6aUqgSGIFIdMN1uGnpqMXxAyHXJBob1MN8maTjiyCkqzDyw7LQCIZi+d6oqtLp
Mar/nC7NdkgoUkTk81fnpxiQwrnHlnY5QEmEYTd1+fb4iWqeH3xO0XPknnvu7zMN
PH5+YXv98hAQHNc7RCv+sCr1k2l6FmpnojhaaXbmRtgmJdvn1BetPvDjNoBDPXY2
Xvk6RJdOqy8YBMcgNDuRq7GLKnX9hyxP+I8LnekNWyFQTWjOqSkImURMyvstzMsR
be9tDx/t4SGis2LEBPWBWsMik+zDWtUqNsf5WQaFu3efoSt3j/ViVu6vsJMQt0t4
dxGGMJU42C1JyeUVEbJ5Bx1TrZNvDHYMlQjzxD9rLVXVWbMPeOXK3sPn+GZElsfC
e1tUbPlzw9VRyJQr0ZsCtvV5hz2oyfs79Nqwkj/oWtA0lfAdeDeAKiK8wWL44Ljz
H0rxLvenuy55XL4xHztmuQQ41HFyCKIOAR4+GZOSQ96hOqZGxqeIH0zjthN9uXtv
6WX4nKGMCp/zxO98IuWbnyvJG0VC68Rx/vieVCD9ZTQVjX4jgt3JyxbapZineSBV
Hrz+7Dg006/kSQC6iwtgupVkhtO7boE4MvIztCDQ5I1o08hiQE8eKiBnuZPOe1o+
2UwRpU1NUpO/BzjkcbkYB6ck9arUk179Mcq9u2Gu+//U0eqFYUHep1ne+U46pCfP
fDPZO+VU8xwFK8/s57vX+WioKJWz05+cZ2hgEo8cPivhjIOfCDXHuWr+PakfJu3M
8cXJPT1iE8iPUvTHB3Bv0+MDakRzYUoGgUyt39GyO6XyQnc0iewtlaQHDPumSctx
XtZU7T/CkcI+7m1aWuFak/lgcqG9mMNFuv9ijewoyZpPSYkqOAn5j7Jv3eDpRqtF
6hiilNbSg1azowdpK/RMK+3rZ2kEbzJmJwUxFS+ll4cEXaJvjlpLVaGiRH57BFdR
eodYyPkHCz8GbIUJSpzIiJzkHLkobnH0LCNY1pcqvQedTJV+Rno9cFqhLltez908
CUsJyeVBqmUJKXlOgbkewQYOCouI2k7gH1c7Oa2owPnkKUStUppJg7U8VmCuI9I/
JaR33nmxnyPKzoVO1ZQiLIMB5XsXKxBlfwRq3pIcIm0t25ZK7TSKArvoyMi6IuTt
8I6n4Pw9g0XmiNuah5HmLFCKB3WA/ml6ElQY79Z0BOPapNjIqNqs6/WICX9rgGqM
WVwlpK6iNL0CRbn4han+0acBB/5aqqZNBhDNfqb9uWAQKkxvH+bpYvCc9GxQYkYF
OEIDMyiZVZcRFf8cmVQk8vDEWEe4CrbTDiw1fg1MvO6BEsRln/g1TzPYZWiSN4dI
U6+TgXieltI34FIEqDHpSedm25GB4KCANvhCzoyAk3ZzfJzyQAbdWt8xsheGDjQM
78w9dma+BlfCatzV/GWkcUTJpe3hWjP6Z22HtimWeKrnp+OEgCLBWIJdnh5v6Kkb
/LwXfg5tsFYoyO3Iyh48Gq8O0yDfojDrdKINkWK6VvidGE7yWpcAVvEl0CQMqNVa
iij/I38OJ/TLrAVDwg5XOdpWMcosBg2eU/mj3/WctHK5eAC/tllv4afSK3kzBkgS
8MrQjizA13N0hFnWV3zXwhSjbqOgSvpUtY2khQ86KKues2yW29VtmIA9wk/mXUTl
HX3AUamI4pG7ptTBVjXaj2prrkLrMV+RRiipO0KprU/B0FYWCaj6zZN33c80Fs/r
IIIv2AumN/4yOU4bJHGsFjmIUUd36tk1rJCluFyU0Enlxj6UclxZXKCbau1W0O6M
PlbMixI+//3uNWAT7pEwOpXTH73l/myN04npgkXdL9hTL5Y8pZXX+dsLvoTM43Kl
Ryrsuwe/EKLAcoLmz8Bjr8tsR6PbntSCKbZVEHjP/J9RepMu32sWAirREfONs5Xe
7uDFkXTxhfTS86fb9fbOLAaJmx9OGFhWpgZAiTm32igP2ZUFFFfJqU/nGuIbQUSK
LzifFvXYfgYCP55xl9UkX3bqO09qyIWDmX6oHvmiI4HYsUvSTl2oZOdzIMVk2JmF
0Zy4dF1hG4IP1XhNAC7NxLR7sme/oYg2R06631Ak1SKfGC9C713ovbnixQTKhei7
uSfx4upuAGzpxBBRQPdcfEGwamIFkjtOXG8rpXlYx10d5bPxrfTcaeWGlDKZ5HbX
q4DvnyUTsTvUuLM1DMSObL0kHEHUMmnZlBKQOB3X26eHqjkWvqFouf/w+ECMrpyW
vizJezrDkgHl7wN5Er+H8aAua9HZCZ04altVicxbUpOZhQIB7mY9oIqpHA+EfVvv
t2zYDP9cne4M0VL9BfppgZRAk2q8DPQLz3rrqSEPreHC2OsoD97ov9vU3GNcrTgh
RuuqWt7DNwd8TzL3ZZ+Z5yVbuVux3L/qBHyyFOgFLuKCjb5wAOOzabwvY2MlNe5L
s5SudViHVIGmQmmOfPcnIg5kyCg/F8oQlBAjiEG9jtZwyNfvHbamBcw9GlGELEbE
uQeG0eU5ifUwxQA6QfoJuZ3zTzAMfMxTy8hCHKk+1pBFYHwDQAaSy5eQ4YuOJrqk
CF8PgZNADSGwLDzEguIG2tr6E8RMbsRCf2jZduHYn/PNfxZy33dXEn/HYwsitG+/
PgupcGsgRNydXloKkCURJQD486BJQag+PYSzywT2DkbgdmOYTClaLqBBwuJasXx2
8YLMT3epcENk3jkRfIO+pDGMYRbaJ1WO0K9puKjcuTrEUUrF8Hlrxnx4+fPk5gm3
+AgGnXtl5zey5AksoCdyGde0uvMeW4+zl4gCNx8Iqv1N8t958u8/99e0CCzN32mR
iMcM9Y7flDQDoZ8LXTFzJqHAL4jK3RjuN0AoGLnNCX7XwQkUlPXRVN71y18hMQDF
1wn2c4XsAuEF2xT9a5066FPhaSYa94fbCzNO7l9Emo+SN8eeZulzMvPDjmumFy8V
qkkC7eHXLPM0xNzgwQtuA6k5jcEwCrkPBwBaFFQzBJmbmll0Vd4wl7LYsYcJZ887
B7vzqRmi2D4oql2v4dtAq1D7eT5pDbksWAtqOZysLiu+JJo9wxSlR560qeT5VkS5
Iyxtsre2JrzeLGSyWpQMGRa2i4dO70kD2g1uZFmJF9+dpwnjNpcpDVlOn0grKzp7
pgkG01EYN9qMmTEN11h/KzyNLjmfwlFEpU2M/BkluI9vuyP6vz267VvGzPgC8oJn
dr1UCFkxHolaenPs/G2yg+ROJVa56+sgnJvnF9johcFCF1/NCdfMXIgh+0R/IcQ6
rTgndtpEI/hHpBASjCxQMBSppIfLWdv7VO2qUxSP5LAr09UWwl+Nf1zTBawQx1pG
ZVo+jDhgFwvTrnqTIZidrNUY4VP8H5eodE62wU57kcdOwanyRdWl/5kdhtKbhmkN
mLZ/5B9C9DBbUC1TJUnJ3I30gn3x9AbnYNyviG0QW9OliEUv7u7HBJk86RTfH8YL
7Ml2zS3QBfiWOiwv02qYHOBXlWYaSpZ7tRTgSltgsgPafXWCIHbG0c6pVIJ6Ng4M
wafbW8UMD3rLttXvKhdV9QrMaV2ntw7XK4aMQUKj40KQSBtkq4tlrZnbWtlh+aVd
AARhxaEO/84nJ7VmVoDGkwhX45niS1AOSLL89zBKwqnfLOnSfNCya0+ema97sxYA
NtfwadQgyaV6pya5TpM33i1kgL9tHSC/9+sKYYADlq1l33stoTRfFk6pG8vsX8xd
fR+M1b7I7JJiZ3MUtbx4ZrTe5dvfhGLiLkQxktp3SDa3EMpPos5As6IFPd2o3zr3
pg+kOjfBnFYAkHVmCyjL5NxGdbXuy68Gf/sruUZfQds11RNdnQvtLkpkiX/uyg/n
lxXrP3taDYV3mkPNIbmiWNTd9mp0asolYNNtPCoAZBTDsvqdiZYayWr9SPbZ9mO/
Uz8lOb9duWVq5hhxquQIvxHhzLGoA+p7y1pBgsGjdhsTbU/AhkC+MjfVU6fJr2Jl
HYRVPCl8YdJrwOdIARQ/OxeZPVeoHT7E63PHdza1iQ6BXWkIf2chFw7OwM7j/9kP
ca6hIod12xjdiCmoRHF1Qo4nKRIWHVRY30PPPB+82tGluZWEuasIddUJraZ68dls
K2gtTpcQsnKx+iLz9sqmDG644sIiqsWAGnTVhhI6v0EZU/Dz6i46PHIHcY3z5oJx
FFcD69rGOtUU6VVVzMvfyTMFFYcrE85SDgj61ch8VwgTBBYOb2pCQ47zTrGzH6MG
l6R24HL0PWiwyv8GCdxvJVaz3B7xgqotSu60S9E8r3D3BKFT6tw4vUpgv86lf4s1
VrBl6OAgXrSLFSOKiRvrV6C4yPJlhMcBSrbmIru5LBcfuEFGyBAWPXtJBYBETVrv
lHZ61U2I59vkIlob/3hAhIjO3wspD8VQjV7oeqjQnvj71WvTQbHZL1PwciR2JsA+
REcWC3ocn1PqWlKldfJCIQ6u37pZ1CZuh8s1IbNDdSBOPu+Nd86dBSajE7Czeb0b
lM4bCr9P/jgHL2HVf7DVEK2IC+iTKVQ6Cwr/jIoNcqkAQ9BqdMNlAmCQbf4qJiN1
0kY0fTwzRafaBWo6J62YcGJiFn5q1Y/vULnqjkH/jsdIGGItQVfmi/GuxPbsw62x
QNBp4KfRGo82xaIdhrFr235aYYP1FaJYRYxfW2wppwObnKuihWvKJqZyhpcA8GZO
TQVyhddYbQ3pvO1ck/lFt+DcXRtmiiTjnzSiiO7Dl9zFCM4xmoCcLv4yxzMbOXFI
9NrBrHWmZGM/E0CeKeBao4hBjy7skk3RQYtiyA+n4i0eDZ/cPmy3GkPKar1ReitS
duYJ2456Aizp9wxw5PeOfQHHd7efv+6U2fIR/K59cNLm2PLWjGZPaScJy1Ab401A
ZLaSRn5LGw+QlJut2YhzxUxMzyD0o0lnHXFyqmCFv5e+2aDLPh88kzFu1Ar5pYYd
eYLc6FH01CKw4GnTJ9+x0fiWw3x08YbfN/Cy8xNhS2H46/xSIqLEp7VC1QlziB5z
i133S3pmihu2j7GIVS6hF4s2egaY/Vtc57+6tYn7rlj4xSx9HdfA8KoSvcKtU1Ra
csKKCcZbJ0yh34NvyMlx0GSJ+xI3zmaxyV61RS58CBm8XBFP5T0naYejRbLe+DP8
nv8fdnygUeRN3LcWskou1xprT2to0ffpLkVLquVLYId8tVDTrB+5g+PTQ4dudh3T
48wG01Y4lTKsQy1tCRwuvU3rY887PecTdfrSxzU5fXXDGAprylIGaUXDTHJBgulQ
87rNnfC8dCbiO+sa4DNYBzLz0okII6xEA8GRJZizJxhhb5KlzEHJtMfhHo4g+wl3
tyU/YPPAYex9E3UPID8KSmtVZwSt5DOL9TrCpgMHtDRzGEvArt3urU75UIdtZoGz
l/uDx/r53rHyH/iHuU4I65YFKWt87PDUymry3Bql/ltytMKsYrzipkbZQlhk+Wlu
5S9wW6ktDxyKz9Jo7ap4FLHvcFmCMpqjpwIjCaVW21pnxK9baHK742W135Ug1CqS
mYWUdZ2idoBepvYb6w+jKnAa0VxDBrzXf7OHtEM38fw0djcdGmLBHWjwTWS2Ynh1
rkRwpr/MDp3l7oNrShBlXJVTFTzAoM880tu7c868sertfJyle9HRv5nMPWgDXhga
ZGMTrbJvFBjsX5zJDAWmQixk4olGG/7KBoB6iNtp0q0pPBGeBZCph+JpQn88BrxL
vqXzS1euf4xWkVm+490AN3hlIU+rbVpZbQ9PpVJHCGCvI7g2SEeBM5OPUhdAviCk
giUUFf5viYv/M2Od8sXh9kOgyMtystBBlNtYJl6Nu3rjyxu0DwwIRRmdNDjhtZWt
P2c2oQm4SWA5/lUAVpGEO7URVIRROZDN9fI+IwAUr6uXichE07RN1rBUbNqprEMX
jbw/CqkpJx7oapVGP2iOW49Tv18/N0rxQ2EYUy/dQs7m8wnFr4TAcEMW+YsderSL
q1kABB8syaJFLYVb9gRTaZdIY1xydc/dCmGeLsnL+WAyk9+lQIFpaOXemAXUdO05
JB9xqSg30m+DppeSIEaclHNm8fmZLkEWlvPARA9yWg8aCu2fA+4/9U68k5OjbZK5
U1GCm6kdhY/lPm0nxrETjbW5F8FTvLnkpmwYhiwawrR+E1t2HPOaASwbdzRgI1m2
EZTkKMtXnKl2C+94i0c7XqcKZy2v8eEKzDdM+LgiSphrp7v8aVJYNDqPhoie1rjD
Ci4iHWv4Vp1HjDP7eMpMvdHFF0G7CNjxip4Tyr9jvu7Sdbz+wdDkdsXABS8MxhcB
Ho7N+pvaoFTidY6c5kawZuo30pFkfS5Cji88GIeCYez4T1KpJRhfMk/kXvhmI701
DxJKV2AutUQjbUN284MlPhxCdCBIEJ5jybnssPpiLAxCF0RPRfd9Ivckycgnl9Mx
FVkSoZ2cRVLhMjTkTdJJCRBMm8g00MZRZ2Qlum9XX1Ythf05pTENWVGocYcqXA+s
oXhWn1b+ZkNmDpo82NpESzb+sB+WAaLcrYn9DQ2DuEIN/tqj1FDg0CcRvVInyaud
QY1LLYYWbOoHbWtp0U86cyFzjU9V1PBwJ+Qi2Xt3KVrEXlrViPk2ij7bU+Qvg1PL
gukfjABrP4WQg684eOwKWwD8HLwTQSIuUvIIesIiVqmTFt49Z+Z+iW71kedxK1Fe
n7kWCTCR1D+JQVDoRI6DF0tOp0oIWmJ4lsQnbFHWiGmNkSxjWkhN9E6zqat9KV6E
iDtY2e5NWaoRIyadGKWCJI9LnZA29kvi/NBmS+RTvBdOaboeR9B2FU9flUdq/OcI
9IEHGnXx3vtsrIzaod4t1jO9q/EXxkz4BMC4TkSEK8eUTdF4YHe8Byi73SM5J1sN
mWt9sfZvVVMKZkxKGUO3dpsPNdgwXjwg/NCIIaCoEb8lcE1QKV/fBb/+Cl7eQjvG
6MezJ1OqNfZXkqWG7YQSlPGcJ/MfMJpxQW9t+OcoyJEX9bgkXfIgRTL1fFspJM/d
uM/twp6YX7IR34tw0gcaKYXVYbDw2twXjDLiQdwQlmPtQY/0kZFoHfbte9JYcr2K
VIrWm1fyN2pQylwukHUKMX7MFDImYhm2eRgVpHR8348/v3mPeLw4KQ+fCb2BAqKZ
5aV5Yh3DoXbFhbn4Xwy1LwI8BBs4Rr2XyoYq2Sw8A6kfmFX1+coQFYLHMHaFKbWj
K/V5NeAoHl+kBJlVqYa6dnxauMBjl4kNoh/nSDAy6bdPqXb6FQBcLOsNUpWF5jon
BLr/tUccnWWX3Weyvj+3SCDNfrPIOm13vyY1ItJUmAaKGNqTp7xymfMrDgP6wZXs
EuBynwRNmPaR7anEcHkqwHECNuz0qfSV1fgAD/6Bcuaio2LFBT56QoH1NDZ7vIIh
qpBVTOf2FwnrVaLCq5CU22ansZimZkJl+5XVd2egCs3t8740WI9m45uPtftyrb6/
Ue1tQO/jV4JqtTf1y9K1q825WFdE76SNUyIeQqI8HozmZzB1JsWIGzzXtvEKdl6+
cXumVCwbniyFgL46OIFMD7YwQkCJbS2N5+rsB1uOvGouBVSNM69WjGoMZK16yMyh
AsyIKdBSSTUHbzecYnj29hK0x9P5Jtf4WTQcpBzdD8tGndCy5y2fgjn2PB1qzOXk
yMc0CE920GUDOs7OdBNczhP2aDnDeOZUhC6VpGbb7753iqP1QandCpPjHaTcSbOW
gFxs7GK5VslffAVu8kXS8WFWnk9KJEYPf8fGJrgIZxTpFTtUVoNdcXOHx9mckSwp
bj/xo/uas5oH8YnN3mA66YxaNSWgDWM+rMkeHdCw+IRR3g7be73vW84AQ8+QxqUV
MWupG/yoZivu7+ME06tkRCsNPfV7/I3ToIenSTbyjIWE7/BiNcO7SYkymaCpKht7
bXMPCHQYftUgNV1StOI9v4wWAGyoKBmlFz28fl5XJgkQhCcfYewoxhwalWov7L+i
GGggWphE9f2bWM448y5qcN1C7LluwQcRxI7nNxUWDOdNuN+NJZenMC9iNkcUZuXN
Qssa/FeB7gwem+v0ktP/MSS6xC8okNoTF4Ukwr5ynSBUC4KMX2muOglt8ZB92HWX
3d9/UEnTW2d1Z+cQXWyOCj79Y8KCGzA45H4+VS4oWq7p4muatyr4545MWEmjhDSj
Z0+ycXsczbbYLVzeCh0XnwGHBgRJEBR4WdEgMB2X2L4zFijYfWHe6lyH4uK9v4a1
GgzQ7rDH0Xstw6TubeQKQOJZTueoDXn+CrQF+EZZ4To4DaNpfI7tALvtadHrWy0L
4g/PgwGDdQ8pspBi+rpblnU1rP+CpAdA4yR5e7SG1wKnLaoEO5VIe07kwYC2TUhu
tYFieYgcuq9aUD6jmqZV4sAAR6igPLMKyUnBRDvhcPHGD9PNJdH+Im5JINtLHNX3
jVawTJxnh9NJ5jU5rd/FPjVfVWsdPuuYq8meeW42PUH7xS/CYgVAqnskakjg9zhe
WY1IRi6zsmzSR/C6sa1beDDOvDXtmID/M52QrQGWcR13uR57ds9hWvIwPJNgA1mv
L1LmIQqUoIuvuHfouyZcUDuU+gAC9aaMJ2Jsbx6Hn0K+9ncw/ESyRgeK9EYLc9rz
/ymC/ixftAof0UdiX/XqQ/TD3bvj1I6AQhGJlKgh2pHLrFuWWmdkQm7yg3zM6lWe
EmqeAMyNg4A4AgOqdyten+6HKGo3PpqZgMVcwBdCDaz/fyJnGa+jMA9jlSr8SE2u
21RV1N5t/UN5WDXJ6ZUGpn+prCQdGpy2tjeHOHYb1CRXZSuST0ccQEhHWbq1+H5J
ZMcq1OeR2HcOb4Pc41SXL6QmTvQFAsG/Jlq9V/d9fSqAhP4JT6Z455DnjTeEcfTW
9vLV+fwosl7h+duQMq3KLNm48DTUjwFEGD4FJe2VCr51epdPqzyCCYN5Z0VASuaG
/UQn9R12fqQF46RNTe3fL641Ggode2FB6ZIE0SRrCfnhxfkl6MXWkqkSDtEaZd/N
Ai/dAY9TvA5jJjdL3dug4HECIAeJ2lYbiGObIRh47NZJvj1WBgLcBVBCGTPc3dYf
bdNkN9QkQTUJb2U192LphMr6j+AqGOs7rBMxFOKrsSxMLnEqKXHVmM6pIzGK8kRD
THaO22LnaeEg4MXNSpwczbLJ4Pzv055mAffuHlJMVzxCrqoyIisPRF55D2c+YQdE
RbwmBzKOZNJwIFgrTJAC3Mby5sJpUIZAOm/lNpoJjk+q3ig79F/eJDcob/ipntCG
C5feKqRlDFG46/0IjIELS/Ai8612dt656MeFY7mS/RSXOmcpl8/0Gl2XpKsUUqmM
YLePv3nf3iopERHkp1yOMFFgGfM0B4xVvArirWEKyl1crXYOyzzGgs2mCbtNFKWK
/BQoKCjf55INSZyfDSJ7vn10QhiabiQ39KPIsgjLAR/ya4WmedUQuZ7M6fd3tOmS
cIja48TEtbkDdJxb2Jh206Ml/dZDDOVxPz8H8zp+S2/698GzzvXfur/2YnZxEYBn
r3/ABfZ8Etd50lD4vpjicHE0O3HhqI5SiFZ+ZesBDO0TJjWQ5SzsqPsKIFcN+ZJE
FLWnjNhheFEr7/QPAfOzUTgsjRUtn/BdyO1US2AYPcdx6jC5kjyKOpwYZggNuygD
dFlsBw3JiZEz4sBXmSinxXYeVvGLEE3hxPgyHm4CBn44yX0HihhET5ztLf3w/5jC
hU48XGPyunLIUQA+wuf6E5KJzBSB2+ab5IbiL9ZHedRKYEWAaK3t3VIWWELfMRya
jcrUYkC/d1p84BwVS+HhVmehe9cZIu50fyqI4aIxw+jVpFC0mxADA+MJny82Vq9C
iMEvhSa0z6KGA1OvFYG/gNAh0KzBrSx7cNDbnrlURWO1FcNmkNPIHJeppcuT2+53
syeM+Syf+YybwBbAvWc1q7KUto0wg9nD37QwtT4ZBSOJVdFmk9AL8H+/SVGYjQ+W
Tp6W2NPhfmHxM/TX1Y4Osw9anoSqh+tLQCpfpiLt2etvyb9EKhpINhR2ASjaA56M
xbMeaRorkv+LhemtIrAANtqNmH+Jd+6abyFRVfoySalSz1qwUdCd4lU9wjwuq9qv
+zPJyePhhZ6ziJQeaG1jMuK2f++/yW0E8yFVZSQAfmlnwr7QFSCve9etTzX7AReK
fm9TeHoCKGQhvjl16vxZNf+s8BD1NA+2rQMFcsQLntH8I8wU60OTr4TERB4UZWzT
UwWKUz2tc3Lc6V214BO7aoIbDcS75391XvzWRscaZ14GYImyMJpE2Pm+ykfAXwOZ
WFBnaqnxvgiNwTu5+kKWUGcbyvVfMNsGdt1DF/PyDQwW006yYSV09vLrC+JKOPQU
zQIi8bMMWN5HPy+f4cqY10e3nwyYjq1qZy6FrJrE43jy9ScjCqvksN0+8Wy5ECSa
wc4+7iGATjrn1M8h7oYygV010FoeaH1302a2wk3l6LV6afJbzJxwwWNg/orrYqp5
bKJiB0d8TxyILNtJoyf47ELH1/2ArJzQpp46YuP/vpiAtuKbJo5ck+MGzMp60Mmd
864ADgIQuu7d0j8a9y5UG7qH87py8oF5Lbj1BfLFG1CziGjMD64h3H/oWV7y8okd
M+wb7231K+47qMltAVgHu+GimakJjIFoe47iweWhCLCb7TWzmKbn7ejfD1yzjDFJ
PtpP3K/w/AmowmodqM3wB0OiobMtAnKpU8MM3N4o5XlzMWLm/S97pmlWdsFjbF7S
5Uc9qGnV95uBH+MgOMpPVvt+kUEcnqQC5Hcjdw9ru4EmibfQ16agsGbVP3Vz+r3A
mmDCptcP8ggdCKbrQ/sdjShR4jkum0IiZGflQa34JKcreHs9+kUBfvvwUxsV0xke
VFDWmFsAXIDg+4hgWSZSeb+hLF5VDA50JvzUMmsBPzXZ6/jJOBQrpnHDLeATAw8N
bp/5Yl/m2jp4Pber4fn64YFst3ulCg04mGVRd3AL1KYmlxnjBYqkocyWflBU+U4u
t+ThumS6V49SvJdOww1hdaO6HvmTP4qeUTSEO8lDBLBD4pc0qWmYW3OfWkpQckKk
i6PzbGNSdDtq6wXbZ2O2sbuFfcbf5zSURIGb2bRe1tfbc6K13dPKY0ChAVo1+3tN
h5rXAnOeo7ouknoGlnxNcXk1XXLc/Oh5xFFbniiJhtSF2uznZMU/7lUUYfbLKY+v
c2BgL67Sl+3gCNNjA5hT23O2SHdFRV2HOERv12PBhVIbgOA54HhNDYpJCZT8FzSm
i1iIb4hlTtWY3C8CDwJw00a3+2aZy6UNpYU9iX+6AxTAWLpx0zO7UOGe3scafpTZ
vrr/+f+dsNXc0Ot9Ky2katpDMnct5EOzaPFFrZXO4Lj665IVlRHSHxuRrKxOZAt5
dVbOlMZ8/+Wc+wSWWBd6iRC19lL2GSqu5LVVD4D2cdf0ho13JyRjkzyQmrSf25Nx
CQLQLS+bsWkuUAVmo0mzYC7Va+xWthDgWjXrQyjDzyfsjE9IYUOrhDXclxqz1mpl
Rj4QcWDxK8zX6ui4asKS1zK63ti8LGHDevypIo9/3xCXjARmEriX3ZXSbSli1c7M
HW/li9isK9veqVl0pat+tDNUla9AYjP0o7a9H5eaYUZvFET0sTFsJvAK82wffVTP
8R06ubLbr+BmSfJDv5I07NoF9fo+XjDHGCsi5NhcenU57F58KGInkLdCjPI9CMpC
7MZ9SuaVhPLWwsGL0I1DT/oab15nWFYmVQ1ZFjBHgmN6h0jbVF+eYVLBKDm0vYPe
JFRaKemikFSJq4kZ2Y6ZL7A3zyvjrZDU0Nd8/XVq5P9HKFkRvutWnPO7ryNHKuMa
FrwY6DxBuUCiGf22zheCEs9+HYEJ85X48KtdZCz05Q3pVFP+BoIJ08edv9osltPE
CLyGomRHc/sL3dg1/kXSn76YPtlND/fkoq10aDrbIXMxWLQWlnpg5SwtN2ChBqpV
4Cadtqg65sKXY0pUNsS9+9ZDTP9vos2G5F+mAc3hEFnBaEMiMXSstba7//FeRXUW
efU6IONGPJ2FyUt1NEfQf1bO6EBnzBiSbTOjRFiilGdv/Y4/dXzgGtU4+x2xx3ee
gjCyJlkUESi1w7II4nEtSbdoznx0BOBkfEciXXIn4MOwwuQQW2ulQsrTlCuMrOLF
OZRyWvCm/bfbJcArF2ztYtOU2gtv+jtrPKnOwVdf21+is7XBcdyYbcgkoBnczGmV
D8Lg/aQheJol1768f6khiPTXgN0Eiqipzoxmj7tiZk/dx8Qa+NGvIXsvvXW+tVPj
zUCEhllapPPZj6fMNsCZGn4uhP/i1Hm5NcsDEhJix4trT+2zLXsFkpzZ649YSZ/z
ZklZAGBSNiiHGTlLEkuwyXBaepjsb493lG2OdfzZolWmv5c3cMc1QxpAZN3KypSe
So3oLPNNPbj4i/EmMXu9rojy26hciEOQYx1ix3hrN0q6zOsEMoVo7eXaUVzcvlfR
FVgtDIQVL2+2Pl65SK0YuRsSy/w0BPhwsVZn+ipyzeNqE4PhtDr+eCS7JmKnCypc
/yTl0bL24BqHXT2cYfTH1VkUq9p8NYzkV0lQgBU5m6gR4np+7GXfns+8Hle9SARW
D/4tUhtFRZiD9cnokvwE46FCVYnaI7yl975NwrOABscsKm9KFB7NfPzVZxYVtWjh
dfwCvWwj/ef+1aTYZuL7szyzbwp2Fgf5N/1hV9v+otcJT+lFK64Snd7/gug75b1H
hLxNqWKaldHIpaQzZgCct7twOyTE13eOXulWb90YWN6qlMh1CGdi+nVwEsQ3DK0n
RKnIOv6z1ARV+WXghsDmKGpntl+EpZD6FdgyowAarEhX3PHy/wScFgzWGz5HOZEw
TX64kjieQo07j7KUzeQIm54yYUClQn8Z4qx6+DOphl7fy03lMS5Pl8ehb3GX42uV
LoN4F2FSbkuXLrEpB0KvyFFNU3eZPnUp/BEznnazl5yuJIiVRTRg90HkwyYijRVy
7mACHVLuzzhFkdBxPPcjWJV8awban+rHNPqB6WAGW5fbDVnn8GDE1+guWRljL73g
BfcnUXQe4JapCXAZ0HBf1aKfzXCQON2zqA6sRwCvXbFv7j72FvByYy69IWs4vg+u
D4TOiScXWm2kM7/Vcimwiur1AY20xsQ/EUyBFzxvoHRVq6kaa2yvX2mh0ofJzEUU
bQ59/IeekQz4Erkg/W1vxrVpJQt7pe3Ixt9n/4gObwnrejyrjkj697CEJn1lpacn
xXM/oMF9qYiHUkpx0gaPt/dRPk8VQ8opjBnILePsmN39RC66xU65m3ebRdXdmen4
V2dTb4zKsgRntD5/8nayZWs65WKYBx8uHSumEPsCVVhITV8DiiM43+b6sPn03zrP
cufu6RGA2aW+zAkLgzNCN8VRh0l7Rls3KOKS8cWzsYMdbUNAiE8aP5ZHkhwHubu8
KsxQYxLCwZ9SszvE0jW39TFyi2wvmEipQoVR5IE51OiDvL33Ym3xV62utcLqtmeX
paGepUc2DHBMEP6mh2P6S/8sVcXU5ijksteKwNJlZl1ovmllSD+fpD4RcsGZSl2e
SUCD6EaST9GbVSPSbW4euBfskfrQUls5dIpmSY4wWpO5uMX4eYoEA7ppOBqeLsJF
o9JUmRG32dGHwklULnJAeosHpJE4T53IetVoW3qIdsEIrNw7QuyHwGFpzMBaFjSj
kyL+SnK7/AIhF0lFOH6rvbyF6IpNexkiOzs6ZwFViQS7Ge4Ni/ai5zxf088O5kqr
CWSI+qlCHAPpNSz3Hhi2cRLUQVYGKnEGyLxWLK2NV2v/pJEPvE/M0+uvnuKBJtmX
Z/u8wYQ9p4XGg/O2LBtsCaU1dwL63CwBIRjweBSGv6cl32OtKYEYu+bpK40Wm0UV
kDB/8HWTFDA2uJADzvoiZ1vwLwHFEidMzjit7g/NbbQfRmtxk1deOrq5sYjokzDx
sCrefQWYbWe4c5ITZpN7upN29jFdSJZzEOaRmA0DBBIlGPZ0xNESy65bqXcAe+q5
DRCpS4e9224EtLrNGz7pQvG078AW3p421do+q0xDfaVxKxtmjkvCBE+ESEref2Ct
jevv9ZUCVoa8GOHHrbeuG8VLKxB6TBZaPC0X+kM7tXnzL+8rGA01RWnTffPUwMTo
GH0ZCIJhghxfEJ5W11AwfDG0osR3ftkyc0EpiH5cTxSK/YsL+S7SeMtPIwFhduzt
GsmKWsHv5vRPgBTWJKf5rNbCpHvYvPxvxtmrydC+2fv6J4yJfMbTfZmri7VbqqCR
j6bG2rchnhOSlx6M9xNfzONXtnjuVjcMzcBIFJPWlaE9vNM7qCzrHmLK5ikFG6gF
YYThrIpTbZQkmvG0ekYxZovBIc8YrB85KZDUnh8g+mL/G2tgXAQk+5KY1CnfHAqO
Dp5mZetWJRBjwW6xnHH4TLgN1YNmfyN8NhXu6syAzVFGMCnAAyzy32B4+zf/DvbV
JyqIYkEq86ErbEhfcwPqiKuGMrOt+s6caKHXzaJHI9hwwt90IcHi00ayAUwh9xcv
hQ1DRs9cm2F145mkFgWW41h958EaOg3MC+dNi0dsOZYvSz3pARa3BnWmev7/BttU
A9RTBwN2QFXjiECqlePLNKhlGxE+oIBW7ZB0D6S7FZFpDPyKrwWHL4OXm3ErnKmq
vGDAZ2hv8D7GkgriTlKWfbl3gXyMD9f8cO27WOpsP85a1H7rriyyHYS+o91uUjri
7fGkzKuaEujlvkShs/cVeeU8McZS/YyG9slyfFZtxBcmuroxdnMP33/hnkt/zzDp
nOcV4juahaxEa9ekzUqa4mmvYXZy6ugyyBKAo81ytBSY5dqt0sbVwXp4yVdOb4e9
q+R0BLp/LkkwYN7Ns7a6v2powVsy1jOjOTwCoz1NoET6xQtgWkdfRYcbqFwNwt11
42Z7fqmg/4gLMFhpee6nbSva77l5dvN4xVSOAW+Ya5O9BUsJNZv5Atd+t5Svu7DC
Fo4WN9cMbs6yq+xbOxO4rgsaJe0xAnsFoAalZauTiTCPILQQ7nIVzqcYekNINEco
6ObIS4+2YEuASRPLjD3Jq6Ko+a3aUb3N4BjEtD322pRMAPTmdtiSu0qksOYfqCIo
dEY1PtaoutABR5nId4M0Lnwmu1/AJNY6k2R5+3BK8wAVNoicCBfvd+8cySz92Bs5
6FTNateDR/RvWt2/biAcu8174tS9LoOiF6l6SRTx0hlVTqJcKGB1IrNoxzBS/Abe
1T9B03YXqp4ayKh2L1ai3UTfaWjL1Sh9MWwP9tn/ntH16Ll2ausqTaYgWMzlqJtP
PairbVRD16g8RrAryXe+9XU8tsMSEnCyDEtDL9c+iMlN/PeW47D4wVFdTrLNxSLg
2eHIYLFuywLVbNcV7t4mRa/dUfMZNvGV/k/Z+zeJx/fmTzT5u+ytoZcvPgjzfFOK
8tdWT2vAhiijN0Htxa4vceMQtkxPPvx0UNSz7JrodpSB+6Ji7Kh7uKSbbgKZS8GX
rnk6r40qLeFoKx+7eO/s1DR52NL2IXLy9b17fvVME3/yD45mnh2mzd45AL0C/IjL
3K7Hs9uYL5LJacHnEyHdVYjwNJ93NNSCsNDB1y8Ot0uy2EEDMmuyEhsowoBdYcgY
L2nrZD0LktC0wvn6REecGhPkHWTGfW7xdMn/G+ImMOJOXbZMIRd95ALUzzaquE3L
DBfwRl0quikb5lcHw72ICpjr8BLBvsPaORsyJKlVaSdUZoTiwfm/wvPv/bIbK4dD
hCD4tC53O0kXQvGUFnmfKn5pXZxRvf+MycTvUNdEMRA1d874GhlH67yFhtsUdFiQ
A9GRP8t9VxrJrZ1x6Frwwc6XDuR3rb5pslkudNjOTVqIxifObBLWztWe+5jGkok8
75RItOgxt7+SQYiNJ/fxT+c4DKeUS7Wa0q67pg4bgJW4OO8kzCmZIWSturl9xNc/
36BxdeCxRjUuRa3/zF4g8e9bQNabKZcbOyZXBblrDYZarQ/UFC4zxOVw9Yz8pvY6
qDbdt5qlpQVQ2eSzt+DyGikuszwZd5SCk5iZFJR9aGNvRIF692Xq2r0HphL8gOZq
DcqGGblHY/r/nkY10eZZYG0jY3IM1JmLD2tIjhBaHLBJcK4e4mLC0jKyBMAhfIBM
mUlbv3Y0kvbn3ATZl1zDfC6uHGnCKWpEbZsut0cFn+aL6ANLK3Rd4CJ24tN4hqpL
/BjyliVovrvsotJCqBcBIq0y37+V1+MF9ars6sDa23dbI77QQjtt+BhO9ZAPLKe8
qKPcTVOad5aSTVX1wNpVvEFiQX8cHu5chhYwocCz7NhKaTKeUHfrm1AFWqqhpL7g
9yM/n7jTo/5B/HpBmQ4at+8sRd/zP4abFzRg8epzUL24Za6NT1rUS+uTdx5UPOHD
Nwoqa5W6hOQXGHrMd2CDYWt/JL2XMF3AXQJgCEZwpcA1aoDxrS1FkfvUlRkw2oM9
aDRDbwir6s2QUkBkviwqVlDC9YyYanlnbX7iWE+RF/VXqxIX5PbDe3ZvCb9m+r5X
KfYX0P4js+xdDsy3aq2GwgpLPjoPLYNVyrVl/eY++hlluPoZlGlMOK+qk+6PVuv8
Gfs8mNDWLrvIN5xBbaYSh3yLPStAUVPYjjmCSI8qu2qpYhD7rNUJzcB6S/psqpco
CIGk5TCrTB67MjXlUqLSlXgGWCdoEiRILgi7aA/O/rZEyQ7RAOXKeKznqANJyAzw
M0i+4+U9J+Pn3I5FDS/9imxldm54m0rjuiNVmC+QqdqkEZElV436PV115wJu97jN
o20c5FRpBwjZcqoz8HBfykoX/kQgIfS+Cl2MgpEe/RbR0D3FlWbqwcbqPDfOyCGz
d08uARE7eWPbespqKCJOxLBugi5ciCmr2iONCkMwqbq56lXWmjg49S6CKecgzG38
y2iPvVDLPM/RsRjjm0zrwOigeLvQ9rFD9r53e3SnH7cJztaCwfbgmjSy3hJqCyY6
cMYCtUDxO4+abZAaIfJmaKpUOpRnJDRhgGXH/8BuDCXwGwKOIllvQ7QmLMzh+CgE
JQhcRQzEaOptJunLSBUCDjJGclhzMkyc8NSPs5xWm6vfb2qA7LCDwu5atpRGAt+m
gUqtifz5VuXZecDjuUgSOOiyJBcJHbjSSVhJwbuuiV/ZoAZ0HZUwxZ+OZVbIatpy
PTCHRmd/nU8+syiSMH8ZsL+p27TNezTEWMOm/vsI5ct216XMBaGhaBm+15rCNGTJ
IT9VuxzSk9fyUXQ9tJSaJdF19MLk77WPzX9X4HoqGy4FxhXpefA0ERDST+b4KeOc
/fFwhLXN0RUnFPWgpwgMKmRWmeUJTkL+eOmnm0TxFwfcN5BS25535+MioBbn/a6r
+wpWZAUGGjMr5Axxf0CDFsvX2cBH2tGBu23UYuGFlYvVcaQ/GbtvGt8rtyR1NdHt
9WkPMUQYJ+xjb7Gg4gEoDGKWl6LkjleiItAqw2G79/BC8zAdTtBZpIo05SMMEDYj
4Mu/McLgddTc+pXlTzrCoxH0kgR8DlcfV/8grd5rsuejDfO7mFu9ycZGme+cMe1n
/21iQNjZO+BN6i9+Bxocj7KeB6E5xXoD5w9Rh4NLAfF3PafSY/SfoqNOW1USSkKK
JBQtbxucKBUFKp0spAhkvSbbze54Hubs2nWFYm8vMwdDCznkhw5AaJXld6mHq+JT
RsNsr/JPQ3ytNCwntlaJZu1KWlW1Wl8ryAmUXe/IM4d1GjQ+NNvmw4S1ORefHCQQ
9zhEV70Y6EZGMnv8QA6E0Y9/AOMKCygdyDpyjQBpRQCufZkjV7Z1UtsyUkLNs9rQ
et7LC7lxc39Nqe+/PDLdhN0Y/GtWP8bP21DbEPspVej2R0wEXBN4CGvRXE6yNZgx
6zWLHcUbU6IRUIi5Mox3doZg9lYel2EvNK5kc5gxqTasEINUifstw+B3CwHp3hmT
wOcCTF+xxzKHULUlcZtsChjdNUJhkior+988724fo0D1tNdXyDADiRt2D44htiYC
FSefAYoZbj+/ZvuoGzGsyEfBaSJPB3im7h6x9FDEEt1AreuVZyrgsNf37CW5DH3F
3+iFjpw1KeOD268idHHVsp0hp/ToJZ6U7cpZapisCk+9kmRo8BFZ2xsAouHX76Xm
GxZxoGhpyye+VF1r48+yBJZvcfMW0U7yb7gTXOO0YvI9KyQn6McpVgD9WbUOcCvL
OL7J0Mw96DdZToPoJWJbVmkKnfSFv3UWEHaSdGNQeVwTAfLcfN09P1J01MV5f3FY
o7wgrq7v8Na8sEebMdsQfpz8L9DewBhQ0Uj0MWUOgXh8BHY35stGs/OmpRN9HBg0
115Jev5ozgbh+un8rtJB4QPCeBofDJK2z8WTkMNHuO229cwrTa4mhdUYc7a1IHcm
uu63NRsamu+yPlI+BVMsUCwarzSSxbUsEJcH5fzOjq1XeNibvOklDksOsAue6207
I4ehfO6uVF9vGKMHuQMqH8EKw3Qbf3443SJm+VINj/s/sAB9pAAHawPdeGbSIIcn
EWi8lvpY8jjAt6HQjh6le8X9FVu0IcZE4PahFZR7Y/3hlSd3NQ5UzPT35jYIfEyk
igISYtxP488Fc5vLXr9JJ0apySaMXM7mZCI9t4qCilux8xCx0hHWZ/M4r+runTqK
suSCm5x6P6amvzTzjvoWkLWU6AxA5SAzcZnAClYohyrh5vgwqhe56pcbMq5BKU+x
Ita2z/IROxzMDsp9oiEdqgd4S1J80JewyHplKNS9f6rIOadupogFLwbTGqVyHUAQ
WGJggK7e1CMzfORsh7jxofuRNFJ3w9XUg9k/dvpI7xENZ87ugKsky6UQHLlaqhP8
3bTeV1jKIKmt6LmT+AD8E0Rd6dAzIc43WUB7HS+xHxAOmSUghg+IxxqWf0M9/vqH
Tp/ZNpo782Wxgo9ksq4pKXFL9J7LuAx24WMKogwsM1VnNcwDxIWhiCJs63ZL7oxh
elw5dcNE58AYzaY2MQ+ykz8YDLrOsatrbyp6fDXcLHwIRdw9mYai+ZkRcLJiG/qQ
OT118ULfm3vaK3JaH2wC8M4fHWBnOftBTF8JNuwx39J8k84KXYJSXFllTezxb9Dt
+r/HSsMZqw5lY9e6GW6Yz5OS41zAs9JgVKmsTtC0OrtCEGAIgjJ0SG90Wr1RBOnq
zB9YX/g2Xsh604TbOnWTPa539tuv+tanGB4C+MR/CtToKOmUsZu0dzF94eH8Jj4j
OafniXg00iW0T9yI7DQ4GN0zPFrVhRsojxrUfo3i6GUHq/sPTSC62gCgAn4yA464
fG52WwayJj9xpIAn8zaPat7uSFKS7oLLF4m0Q0b+Z7Jtt+3LmoXfMd58Sc+DjIDV
JzNwzV8R/3xZXfINOavDakI2WausSNqkvPOkSfXcP5y1rax7RWs6yUQ7T2Omwgn1
9XMwHeiZpvXn2wLYcv/cuLboxNTRkeJrDfsnwXXcqrc9w7rWm18MeL71VTxtQThk
zp4cJnnMNqiRcG0qo4KWUT+4tegiGQ0xCTvkLlVc6v0RxsZ3x0ITxekmtpvXSoNM
JjtMFkxRN29NXb1FTDOuk3cqipePLK0UMvusLQk9R5WbX8d4DWRd+ilpup5GTuNW
OO9vsQoHe0ygRGNXQGDV2M7fcCrNFCiB3pyL7JViVLUivjWlIQ0TDTebbDAlUK4d
bct5Q4dEzSBKUii8n52lkn+7Bd7Lrz0oCwI4OFarVYdLsfC89oEola2mDqdR7tj6
eqIAtorHqOhgSfk5hVm7t2aW/9rqn19wm/JhhSkh/V68lxfWwcAIhfY/s0Ys2Sg1
KS9mTPw+5fCIwgfG7m/TZy1XTqlBBw+vtJB2e41nN34DPx7iF8YcEtnvmOsH9kV4
PxsEBhv46+po2E9g9ep214U2Qpf/LXO7RZeWpJ/b3+QTWd1yBvB/FfjDVTfW30xP
8cSF56sXvbT2dveLs4Vjxx5d0F3SzocoQil/oRhiV46C1pB8n7aEWDPZ99PITHXp
Z05WKHLxPBfucnOF7ykJNDLcffAVriZAEc609Ty/0MqGfwMmS0/hxoivzXvehFrs
COVhFd+B9m9HEtnKn84CRZNU52VFYZTeq4a8O2o/nOagA13WTPweBwbO6C3Uc5Ro
WWIjCFXTPdpMlPUfM69HK7TqUtZGKcpZEGQqzlvujD/CLEieWAiCrk8vZKB6W+Qz
ZWUWmUtDvBHYLPabEHBpS6piqvuXl+hA2sbd1iEEvyq8X35+eYXWttKV3QHaaLUA
LxRiw2IgZPaTq9k0pgeLIfMKh8sUEbXoT9ZTSsumj1DJIZFV4FaPxIYTokw/wP9U
GCjvXiL2CJMCckL149ItVXQE6XCPnkAviCLSrqAI0fBLVueh8J3Ag5UrDsIr5xGl
brBtTBIsQZ5HTO0Ci+oDZVkfCrKAM/yvRpCHQtk5lIcFlcrRwS1NYt7hFM87jg2w
/YXrQUcltsnMjDa3Nb6UkNqkKh4dfsG7+noCYdGDEI208EqQn1taRakx+UHxKHfK
D5PR/+aVlFUh1l47rneXetwSRQU3CHAXW97oCexutyfYLnRG1wCiA0IOJe0ikQe5
B1F70D5O6T66HEhjLXOgfhYxK2Gwwy9iZSB3aZI8Q4EvFBELdjJkEUBgh1z5vIXP
qqbiGaNFzUnE6oShSox0/3nr9d/Opx3fWIUhv0xf6zIY5uVTt+8BFpjralFUamdr
msvAp59xCXNO/5WvxFKNF3JW3jnu1wF9YGmCNDYFkm90kZfFdLoz+IepglkdqqJ+
tWijFER1YVrMf4qLnNNcbDPnQrEU0HJ2rb2N3fRmgWUnCU3F+S3xsC8n3zXsXdIL
FLLegEbMZuC1mnav/mlv12vV3tbVtPuFtx8+8dY83qS1/8BKD2Gzk4KubO0gi9gv
Pa2WG/My9vG7/MG0KFHgLw5pfIeneOGbeCptRtctnOuRfLCipo7po+T1NOsDMQIG
Taw0yFRLAApfgDjazuWK2CkvxIyyUBYYyrXiDa69NfYDmKckXMK4MhGgNTDzN9YL
8yNfiB7YVqlNkN+Q1QS3B1xLhBxM0Aja2qTgs99+Y4jw0Qyq8062LHSMVqKUKFBG
tAYwEcOcRcXy2yznRyxJtWnHUo3t1L1+woZYJMPKO/stRvwCrV50ErQVUuNLPDfd
sPdV0E5RA1V+qZofc2eRbF3lTq6ZTQY4+kYWjjneLW9RGIMX4nZAFnXQaM8TdSa0
ygYZmYlc3qHQlh22z1c49Fhu5EsTsY/eaZT3lnhxgPDjHqdsx0b8asUuziRdU3EY
3Ykz3emK4DX9W9MhvzIDuiyX7AYX1281L07nsdKt8w0QiBQU2/Dwf0kQqOmgQix6
jh1NCjZFgkcS5S0on9AToFOejcnR8TqeT0UfdbOYo0lCd8fKF2oCmEgs9KvHVtcU
IMLNMFB3fkTJmWPnjDH0beCaba5+14Bf6W1+hVUEDt4ps5C8vd2CzgMbcUIpBnEm
uPWHMlvDL0A0+7l4JZ53yDF3IPLAilsJ5+YUh+ICZEzeD7xVELJfgw2jeavL6bN+
23Z58xnwaTQBd+tfDI6oGieh4v3nVqTtIia/8RCV15yJdc0L9UaKdGc3Gg9op24y
l63jnEAmV+lNMp1QqzJiAfhmWFzzszQu5+leo18Sef38V97zZIm4WhhvLRssl+Pn
wYS/VJxclA57aksasStqAHBEh+JAgPDihqYILpPesyPExzndB2AQ8JyRPsZ4bpmZ
1bbuGlC+15cPeO+2XsgGrog2D7z3rLYf91jvj8QKKbqP/sf3901UjMmYePkmxAvJ
2yx0NOLLOiND3OWpVFnhat6teBFKtGqTjiFLeDp+FgpXFwZI8YctvBFVc3oLB+3t
MlXgHNVhPbCU7vPyeUstb4wmQ2XOoIitZ6Tu+vamiz25vjWTG1v4dorfK+rFh5NX
mC7lXABG7sUxsyYj7ujxZrqpOaOvpni0+EFkZAKjdiPmBvOi0lTHN7MkiHivM9ix
E04puGl/Skl7yfSY7evXm1kgRzSxWlWxmWrVHj5hM4pNqTJ1ekIfC5IENmsQBES6
YVU28uIU59UisYx6ZNA1Mdtc8FCHC90HUHcHhf6e6HtDTZOactUHfTpD2x2wNW2H
yMaYUvU5CKq+C3N+IpZrLR1NeeknqGZPZ/QyBBpgraVvU333o9V0Utf5WvRFfxKn
9bg8ThwdJKRQPOJbdwXxchfD8aD8Uj3jMZHLi5RI7C1OMoZT7Nn+g0P0foOB+C+y
VOr0YfKYUm/Mi5tzS4zV+whuQ8wV+d/w+pH18By3RZiIu3gk8Zmcsky4uZuyk06d
Y87Dg2za4wT3eGBNLnwh2bfOVNNe9Mm5zTBSwCokjIxs81Fy+B9m7BtwY5LLhRtY
Smo0NNKEWrOizlR1elhZ6lsm30TtNoGXnaC+QVzky9LMfg+HFCcFMxrRw90p3waC
4hjc5ghjPHxs9i6KvbcFWVOBgN8ISNtr7YIC20r1A9VbhJFN/OfS09prsTmUMcqb
/N8SJ1b8hYTl0sybiNyJQDvkSUwOfTSCol+vQsLPVFqWIKUjBadxuVJ7/zC8IJN3
SUjj7wGLrwJgSlLY6hSl9OFpBTELxGkwQYgU5C+2bd3mLnlbRB/fQDnyyaqgSQ7r
luDFC7rMYq5FUnqbsW8pqXY2HYPITuvmIdI5Sq932RyAWvggRSHEzNKgIdxRL/9o
2NlWsCvl4/7EaSWUb0MgCw80/dXcSLs+NocBI9KV1ZyRFVoR23EV/iMFRplSXKyZ
lQ8rViMLo8Z0h2KvU0nszh1zmJNf0HV8y1MoztaCVd2tHxkvYqKPWE8v2oRz1ADY
sdKj7Bbq9F5/mF3tJES0lntAbOt2WKCX7CMc7n1jFyMPuWeMIe5eW7IvLJJwQYc5
J2t8DnA/fhy1ri08UVjxKUHxhzSptbm+Kr6b2eRJ9NxuCpZGl/wHbjaJgoQr6A+i
IzXUzmCCFf0afqWymjczNLU76fVmoUBugpxIdgluXNdEwiRvNneMI0Gd8p7TQqsS
+6Brk3QKsToUWp7IjmtkBQ14mtU1QofZwBpm1SMrISRSHaiZxmjXrNjQHYHVdDnW
7uRvys178pYBtJ11G4nTHmu9aU+NK7Xvk8S0l96igQ/B871MyYSQmHyuXOZs03Zv
jzwjsRM9GNPBJpkb24kHKtrDJD6EiFpRlkvSRMnujYoOvE/GWg71UVF7YvuGlmlc
TREcxSnUyh663/IBCtjHn3nrmEB/NeRa0pU1NDu4AswQsjzjOPdQ8n+JP+/wdNUz
6JB1QXAf8jggCswilCXa1jL9/i8iDkZtF1mqvyu98I8/mIULc4ZeInGtyGPSRBXA
CaAXzJJ1vyhSPttxR7PYxrbTW3OweuY4eAVHceFEitduwmLpIuLYo6FRNNlqJyDf
LMFbYxJMaQmwZTsx/N8kx71/E0o/0zWGGzW8HGV8OAF4n2tbWeQMgg8Yv4UrvZqc
S5YeiF/uNRtf1Y12yXO10uu9tbkfgmZFZKrTR2YpW97YckE4UnsHtWil+8y1TQo9
nM+8Ec7M+5IHGa4O3nPJle7Q4H11bu69Rt7QUp60Ky2C4fkgwpMD+LDSLxjCLaHb
GckpRK9duKsCnArM0aFHKcwXxOQip8q1rGUPxp641s/zvsS1BFwDOO0VySCt4eIr
DoyHAjZxwCu8i/A79KbYc79FXnWldV+84Kg0bPYL6JY78z0NM7Z++KYvUIGAMg3+
iIDBJshCilADY/MoMcZ1nRQ9mZNhWqBasikM4Nd3b14CUhLRozdz4i2ecSA0h9BV
3HCaPGLnl/ZyEarubcHveU405yTIQZAvkwmDVJnjNtIz6M3pib23HJwQyiWPjggV
AUP4EwxQ2N7DjUKMxddrbRSIQClvfeIAQOBSi4v0jCVlIBBd9LSdRm20skHao/78
JhJeouuG/jHH0XmoFbeh5LJGiPfoxEN24y5o7Cu/KIKEWAb4EqqBkVvgIQBAb+4o
Oo/cEKgZLJG3kHX6qmdnWendKTRTHVCVxi4tl9SDDNWAP70+SnwFU4RWkM2t8Aks
B3UgGzBF/uLlugRz+ktmq/xKweKGuOpquZhIhafcO3xJDXI6Y9VCvinQBtpkPukT
IzDb3zZ9uUQnGLkdXyO92QGcEb9fwdv8CG+i4BNZxLWzeNz51KuEaQ5DExjyclpa
bmN5mzhWWoi4k/agrQTBaHquqLDRyujsGAJ9s/xvk4jbNX+l+o95g9qFGXwL1UUJ
vtqul/f3TAuwA7Nb2L713F/YdvEpJ7mpwtbldrowhH6mUR71QhSGdRjk+WuRf7am
uniBm5cRgAAt0MWToU/I9g4iyo1S8sORI+N0YAgr5EHmjGLZYmwi3FYgJdVYq7HJ
RalL1lvFk274T1A0cbIwGI+vSGLPKScYrq4ZEFGYiz2J52d3nmHBzqe6ta4KhP8P
Su/m6dSAFWBwONXBjrt7HXba8DXQUfm4aQl2b1pfcRkWTu/ihg7UkJDRD1VClfxS
SbCyvcJPv/ggAAjTtKAVZVSwn8Szj8psPE7YjxmCHcP+w3SmVZeOATnzyT6LYhhC
WG6HGSnK8+hL0lFqMlZHwAqW2VQ1LXy4AF4TwSfY9Eg+3pppfF0VXy9I0/TLKM4Q
yIDrHg0iqNT/2Vk3MEcZmSrSqiQF9rFNNNv0KHxCvcI5JEPJwlKVEi85v+SUGt3L
rv9V3e6+oinhiR7z/TFC0fGbkegcM/kiS6Oh6/oUhTMp/1ywQqkWIUny7ElygRTl
/LQ90sAqL8SmzQG3OUlt3lWc+B6kQKk1wV9j/w90VKbP5uO2n12+BIfw6EtPXtox
9VswcXQ0ERfT++RzWsMdwAa1U/TmYr2apuMh+zpFgSNdEqQbXGICyEvynGHr3W4V
XQfQGGI5X0qjvG93U7HcvjAIwp6UFfbM3v1KFkNmZPJbKjX69/BKGX43F0+Evw3J
dxsydOV9DJnPe7vxaWdJ1vjrUAwXcmRWMkuBhnEunqY2L7zedx1Zutl++OT2y/Z1
BdtADjVaRAlbBovbDgznuIh/PapUOzuFkuVHlSFRBQxC5gcEg9lQI+lcXD2U+w+U
D6f4x0njgvKgP3GXOpJdjyt/B9lEPmLXIAodtz9LkuwEtuBNtByKwnz6M+PxnBbB
whlPfILj0brD7m4qAzMNl6rNmRTGPbWOzHf2CQ0DmO2y2R/Yyeh99/X3uSv+/upA
fgWQ0J13XmsYLKgPYcAfDxSkAomzeS9hjNO+wJ+dOz2PI2cxfW3PokXxfLE0f+dn
bEbzgAj905euX0FvYpEoJCoumFDn5tsdYQEWn0bBpUwaXU54VhWHwUcQE81Kv3XA
/qzbF18yeEe6P1XgM8sXhuXodU8+fOAYL/iI5ytQJAWy9vIAD7UvO3V5+fh8tQgQ
1fYCuuMBfoREs33mF8JE6AjnE5ZlItn1Y1EWcmAGfYbYE92UZpu+a6A6JbzL21SN
DPx26E9YKxV5swBvZkme3l4SZcTPSSaOUrlN9GG94gnQ/iOddcIeGps60afYJgLw
366RrK/voXBZHycTm3vZOPaEllzKocusodo/BfY4iBV0H4/6iF1sqwDPhY8GyNSj
mBQVyFiOaE3F5B8rtyXD5iWfB2xlIX9K6blgFaKjFs0rTZqEd3XEygLVYganQ7C+
5nr1H80R6oXJ7XI6CkXXGnQ0MNtTvFKpTpZdiXUYb2q6toSrqGeCBgQU+ADmJ3Zp
6FkTO4BMc9DFs6C4l6aedWWxklxiPxPdmR4WFQ+YfuuI5R7A3rFzh9EPb/9Zz+29
2fOyOJoPEoD8/ir679Vwdy/lQnxYeu+oS6HrfGzSwpA8pjcFY55vhw8PmjS7HRR0
6RFfsZDLhWCx9i3cvFrBiV5Y5eA4KT77+Hi+tYlKhrS9UgGhr6yo6btlTjTxisqS
e/xRbQ3xSUfUm+zAuo8jod2M1ZuQHdF3CQwLQiMX1tHIFNpRK4bUXtLCyvxf1lXo
bGw7oe/Nde3yXHsh9m51LpQPgopKmu3lEftQRdVGAJKPtK9EfSDkD+Fu07mOetg+
uTrl8LRfCsOGRc686eA2eIwm6l8nUj6cb/VMpMuk/JMpD12OCYm6MhmiZiCCf7zh
llAeEm2q9I8ob9g/DqkH92MGfB/zowXiDSq6m9HNt0NKCOZ52eBhX2Ywh7htIqEY
4+mPhM5q0d1VJW2h8fJO4Q9EARESf7QDB/jzk32Xgpfr+hYnoBWXCV0I/cT5arsv
KJ7g6qsJ4fiqs4CO0q4QiZlUgQ/U7koSQP+i8pCMs2IZzFKtuGWoBl/8Bk35+SsP
OAv6z+KwdHkkHrQqfXKDCiNcFTjYzVFf5CFHIQTeA9M3Xe94gCefbQqKPZGH6cWV
SSHFipsnzDQ/t6oVlEGVKHIOPkB+v+zsd1HJTPHdMUovz6vdBQZmrO1EHJHV9WS5
HYb5yNwT8PGvN4NRm53/GxlkckiT+WEOcux0+/SPmHu9Jsc5AboyMkrLvlHJghX2
84n3XTY+9A868RVbrpL72/6hbhGebPsMMTQaVTZyAiuNpQ09h+gQES84q+9xHdrT
0OR7Vorhz/uv3fFdNJjdzYRQXI36BYy0yJe9t2qSnPzsH0V6Z25G0klsPTf1lJUs
ZcsDaDrIiRrpPCY5TjwLV8ClQ1w1GOdkNnwcgqbWivHrpYFvjWo5DLXxFR7jlTKk
xbTyElIVnLtC6S7Tf1zGHOZE2iGZizOmQMVuxOjD0uKT5KIXdZySgJa+8DyyqYGo
pGUVxEb86iaDMGOEBc13z49tyxAGbFQ48w4KSKUhwQhYSUp8GGWqGVYVazgjg1Mi
F5SQmc7PZnivN6uU6N0lhNysKhDIc5NPd4CneBdvcOJJPaHPk5mgc/MdQqGPcNEJ
Cr1DXKGdwtP5zVu5jwqwPJg0UBx9+Aieovw6Jyhz7n+6A1CX2nM6WN/XYnd7W3rW
Xxg9XoA5waRvAngS94grllRVWcPTSkHB2YvhxNHWsGj3ordqdrREq5dkP6uJIlWQ
jo9956/w1pv1UXRadPk05GypuQT/99xj7NdB6K19nR4QvSPZ61Y0VnHHQDszoKQe
GUmQBwDovIvRCk8QaHMGtTvtlw4r7FD1RQ7wUre7ioZAmEG+PCji4RLSw76ZQ3G2
dU4BeR07txTqzmEM2na1IlEYbbQQHZcRngL4JGaZwI0MKi0QE6jKwOM5/4CROWyC
NNsU270n9y1QTk5WAsOlMUKIHxTKvRu0ukdqWeEtpSJPHN3giTzBDTg5ISZPYRXf
dbPX8l3j4N0qiVxHtuWKWA4ep/i2EN2gkgMP3IP4YMy/Ejeu6H+GUR5OF9nPhH3h
nAtiqYrEAdqOqzYRTjf8gNXJKYa51Ka0y9w326S2PVw+CpkDStTv/MACSolawkzp
j7PNsS+IfGyjGwUazKIwJfbpWXWAF24hIKqmdK1QkKW3/NK+jP/WV0bHNCGb4EA1
hjflVvQIC5VnFknjdzedl1OJlLr87gljPOiQsYNxOeI4kBM0kU9BCwggGn8S4MTI
8zvonKd+LcvfRbTUf/26e884K+kKv1x695cQBuFLmbocqDYl4byKbGPjZaNlZVLm
tobf1t7vAZraAn4ydb4FEbmTk2UDEVanJc9uOK4U2Elutr6//mw3VqEX3RpSkKvS
F+dprWzIWWEbidTwW/I1/xkHH4h0+Q/j8Rn2J9a8EK4fGStR7sZutoUzPphikp51
`pragma protect end_protected

`endif // `ifndef _VSL_ADDR_ELECT_SV_


