//----------------------------------------------------------------------
/**
 * @file vf_axi_cfg.sv
 * @brief Defines VF AXI configuration classes.
 */
/*
 * Copyright (C) 2007-2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_CFG_SV_
`define _VF_AXI_CFG_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
VOlbHDfPjq+QuLvL8+hp60b/7EQA3nt9s0jDUK3VV3tf/Sn0tFZW/Pv5wu+uL1vO
dEQXMgwIPlDSuz/Bildc31o4Kcs/jxJpYgAJUYpvezX6EQH8N+p7pbFajhwWsMg+
ggCbhrBdtFzlJTZuoZm1oTdTd3KxpGHSKKdSCrgQmwAmGPpz8ewzD/brbv+u/kAn
ykCRmO1c53Y/pqTFAk/CvlAVWFxHsuThEjKodLgj//rK4G8uy9GS82XttjU0sADC
VEnHfMlyMXETsQdbyr1nbLP0sJInOzlfyAKSUbfprtrPuLEtkbRWKYx5KvGpb20N
1YkFZHOBUs8kS5axVe6SPg==
`pragma protect data_block
ZkU7ZrAW2ZjtDDJDATSRxDm7Kl9LRjUHh1tSGLgRMmXmUFsveUs0GhB08M1VrBzQ
pk6cNuMLa5gyMsSUhQ5VlYiZ0Dqfceqqz69GCIygCkrIZCFUYAG2vfP6a8TTPUXx
M+KmjAafntn0LUY+ANmcsXkHl/hRI75B5QtUCfi5d/7OE0dftxQQEnXPlGzypgPx
uzj32DB9J7IUlgFMLoKiF+zOHzN0ThMWMZ2uT91O11Ibi0+AUyEWTngf2SYjuR2g
v1R4WhwOPFQe/o9oqvfdHv9N2eo5HZxXzjc/Ll+whrKd98nhFymhu090/qAuNnkz
i/9r9TSh/QrYjVHLy92jiLT/21RguI6tbTUQhE6EYCfiBOL+bccV0QHw9cHt9vil
jXEslmHu/uKZP5YuSwG47ncWiDEJtkdkPVypV3qbgbTk/JA8mEy/JBJ4VXBIuTki
/GVX4Gj0MiTWXGFbGfezXYvoL2toBN0RtN0jAyc99QhVYqrooMgGuvVU/qFKIUgg
cI1q3HchKbQgMyIjyk8EGnM6/zc7UaXnHifdSUJV5HTZTxkK69tA75Lr1jvL0Olr
QLj6eic840jkgoXWGBtzy9DgtrOrt/ODFqNXQ4BoV1AMwsxbZpTU5FdUHeYfVaNi
RVyLKMvylWEGQW3HCDaUiAnOevzHMNrq7ZHPABKu0UhP3DJ71qI4/ZWrAIks58vh
eMtB5ucNkqRF3QbjEqwNZa7KPXgUGkWdgzBUz7kYQOKOrpVt85wCqF/pTYFsKf+l
k71Bt2VQIg/oesyHmJt+mWX5DXoFOIRQSB8Paf+ifl9V2AAfsHUmLol5ov/kE4JU
OEn4TpJt/sgyJcQMmCw+DrQVdOV+KuUPYJna7pi7Fl5ZNSkQHo2Eti0dbrSovX34
wfxHO/TRXesk7TLWM10Ntlk2sX7gH/l2OCqWP/wPaKz/ic4h2hEuVXw+XeSmquyS
44EMMNvBmULKseF1kGOMDbMATLWUbEjzqNsMxp/ATv3eSsjBC2qu1GvZnd7czLUR
sqG2y3HiAilJDnSgStJF3Y4cbFt37bS6DXJdGNzlOyrYk5EdnMyDj3IiTj4lPxto
4uArh6ZD79w1ToimC+i1mUF14is3SC2oRgfIrqz4N2xPZsmoaN+5PQD3uJE2CrcD
00YG9WK1rEvgFRsWAj509745voVzPx5qK8OKcS31jiOpxB1RzW1YltgfY41/+Y0D
cIP4WbUxXufSeQpxwmqGwUt/KEI+1C+9D7ufrN79YNAc3xdFhvJXFUjXrBolvbq6
aHGLB6RcnbINlhUqVFDeEfEyzh0qofTXVvQ/ZTk2dlv98pSObwhMc6B6m8TWzYtq
sihe2WQCI0hJzwpAzd8Jb0vbKKf1qR00tX6RzcfgXn8x1Bt7abbv3ppSTdxRHHUD
tlNFnGi6mjTuuU6Rtz2VTkwqgPHwKV3zCYBtkYkifkzftFC7ZvH+WG98kuFHpvhD
VpVLjuE5LvJL9SaxHiCt/asIp+UzI2F4w98Zyh07VA6ikubFP6m0u6vlF2EApRjm
sXlp0l+zztuSsZNe7C8jE6hlHwrk5quGYeoV0CAU6sb8q8QmM9xrLTFT/OGEXxUg
6FsPq/gNea9s229o/C8ItL2Ykvl0YBY2qc3d5xgiLYYqRjoN0g3I2+EwIXGqmCKF
sO6sdXVxSRFFvyv2dl/CU0MvRML8pPRwztQLDAekLVmXhg1c3Y0jkirDY5S9rJXg
frVLl34nHwYziQlWb20hTy+7xWfDAInel5l//E4D3j5jMgnRmmt0Xse1FUXphbtQ
deAU+jr82IWRl/aN6NEjy0ysruOzLsAjPQq7IiCsyccpZTOjm0OabDoB3DMkUfKG
EmqVS2wMgSX9xNHhS1HlfPxKnDixOICxmCsZORc2Yp0EdkXeMcp6jAXs+g7221SP
3zMUMM43imluZ+xXqG0rZWhiWUOHoTw7ViLdvfVGC0r0ZoCfLTgWVEbsqdwe0Ikd
QTryFXGl9gJqeOBqNG+IPa4DjlB7X3RS2e5hypqlQoNUEKiGKpBWxKn2QXXMkBMK
4thhZFcOfXbOloW4dSgt/lzXAZDKg+o9+AohlwqOIe+8BHhRCiyZhXj00JyuSuVW
XvDMtnruiC2LrF9yCdM6CEGaCary9K/Pdat8BmIMDpcwq9Z3hel1NE75h7MNR7xo
uv0gYLI5WqqxDZiXN1EMptYxiIZTLA24e6kjYNqAD8bMHlSIMT2n54VBaG9xeHgh
qQbXFdsUbrPKah0J/twiGOMEGovJrrVnEhsDo4F/z+1ZD5mrVOBt8IPOGCUK+UIZ
U6CtpqMmt33tDmrQyuFjODDojv44YwSJJqe9UKqQ8y5Fs3HfHhvKkAfJ4/ffceOP
7FqmjMS2+y4P6+ZSOS/t+H9A4tENK07IgjiD3rOtUe0QP5Gxprpn2V/bx8ALFcia
wL7BMKclAa6Q/+Qspn1SeyIfNoctlO0jHAFVgGbNDR4OC8y8UETPycgXCEKTvACY
7ewSok6jPIfcu4CYMl4+zLclQ8gT94Qj1l3mt8UpsfW6zMQEqxxKeaH58DaXIBnD
mBnevSoA4OTIbTXckFAkJAMp0XeNoDwAAryCWg3y6hRSgMwJ1CXuqBALuQ55O4V+
CrNSedjexoCBA4ADWS4DpjrRyN90jAAB4d35klw2nL0V+gWfeZkiJ65kasSr+Mxr
bpILNdvhvvC/pQifXN6Jkjrm00DnTj0Ygz2ulumtllPjF+nLOfOVjtW4IS5zRZ0k
3Lwjznw/W0E4cCWOnTwkluuVzmyIXrlyYW9vBvnrhfkboyPJIKnj98d3Y78JMDZl
xf7qAjG5TLX02rLQFo2bVj6ZCkcCu50teNV9jphTQuuAJlJ02khIRhSrlhToJWfM
ADIXJU1wyUb0UWgLP69ohXkcUZfXNCTNdQu0lxnV3bq/Kz33PwPCC7W8ru9R+MmE
hUh506Pq4Xnid6CpkPtrLZTxvX+RVU6Ffqy1h1ZSsPTUYkhM6KUQFLoOm8IQ+0lL
AtU2G4sGbOzEc8G+tZ5kKCX2jdX9VFTuSs2CoZsbDH7n60WunwHuQj+vbXjI+0+r
tlyeBPOpRQx7D6lGQ8t39m1MysomKnhtymSsDdngoo6OSpI6mo+SW4hFzA9GIo+i
wAB6J3ml8JJqaJFlqE6z/+Glae9GySFidXNl+wZRmM+ksyZR+70Ga5Ox2gf6YC1Z
pjnwgFXYuAivi7A275jetXmRmwcFByRI2Bx6XRaMJsQEtFYoAJ1xC9sfkSNKICQ+
bXX2dJeQaWBKjJIbDeJrvwgu6HDcX4UnhiOyZZFJfziQ6ZaZAR5ZOGLeaglHUC14
/TGJEv8mOy7e3NNoCpVTvQUbBNjdWGBI/TVz2f2GZErejyXNE2CjKG4Jyk7K/iD/
LiDU+Qxs+zVx7H+4/R9nv9jFqI+cTzjIS+CVwHm42D0HBW0ax3fTjc9PoooruGN1
X449IrXoAqw6lQZRpklurKgx33jtGHCpOhoovCnFUCxwJsmgRuN6XCCcywKXYv8G
57UEKVBRhWQYlAjWZpyj9/cIwy/rXMXCwtlHqYsC9H9rIiggHM/tfhn/ifEEFzJq
EEdZhiYTnfT4JBcAas343hC9pBYd3trt3X1AZ2l7564Zmvf6a/W4HnDRjAVn0tEc
ng6RqRBrRXmpXcR/JvEN5R7f9p8s59C0ZzF2qJjdxruzfqg7RB6p/bUT7o3AERAN
lbWnSJk76qlXW1Qp3vg5+eRp2npmBbGG3VhyozCRKJAgmMMufUD3JUxmyiiKGNAX
QWGNOpJEYCMtJ5mVh2fDsEQgG1DG1HfxKzc1dNke1OTVm7u5BeYqKkAwVwM/ZJDR
ZggdkpF01wpA+ya/L1/WcdM18nyEtYjdDSHvqm2svGer3WkEusJJm6kTIrj3vfs8
Zw3xrbi3D0u0/+N7qoGg3WzV7kBnznamRHQToNgLjN54UbxaBjGWCElPWVvJPW+A
bJPkSwGYD9LE3/sQUJdnTeCELz7JLcchsgD0chFK5zUrKBO+dKKa/Q7znWqvFdl5
ltnqR8mTmzkzsLUzLyvQSKG+nKkS89MAhx5kUKTRdcJW29/nLRj95RSH9X20gpTH
VTmgZ0gB9lL25W7CHRbWSbfKtarxuGDaM98kad+eGtipDoITte0Ee/ArZuoRJvsU
87P34HF4icUkbaKGcQ2ezL8TVnS+gADjBqjloRgwYrcGQT8YPSZyxu1RaM3spIJX
hPt66/xKnN80t2nHVTfOifJMl8FTqqw83P3DQsFb0qsQ0VXb90jPzD8PU2Yz6Kes
8c6nMBYZ4FOiW+fkTg2D7ccbejW/xvoIeAvpaVlTz+haNczInrsboKPr+4zYizgb
hmRN2kExBkXOHehhOEdRUtbhLWySTnDS9CrYwnpVI6ZaLzceL8EeKKzdefRZL7Yg
AqLq3xEKMAwdqdGCpgFT1ynQNVtDNR49HdWTi585vUXXxuRNmUC7q/07N92/Xlmf
iWMhcHcH8/ZX2YXsq9eyBFditMIzP59hr77foVcgeW5aYfpXg8F6kyBzSBsM3/Jk
fdd3135Kozp6YckZXUxeHbWY8pKYlWKfUzIPhe56UInQmSP/TPHMCvbi2t/rqw7c
wJpc9UY7BY/zCwM1iOLvGUY0O69wZKa8mwaXwM6cYGMgjsK37h8rJSsS1CEQCS8Q
HfE/0iz4i+bPg7jNmVCDeZnh7Tf0CkSKKLeCa8cCNACGWiRkcdF9ULTUlKAnBi3r
+dFcp91ulU1Kx+Ddaf/ZScG/ro4zIv2tt6UV94LqQYwc2wttHoXAVOSjqmmV4pZ7
ElUG4rV23o/eFfpBhZPk6UJy0mnHzB/DiUw48EEqCLJSkfdCCkwbmHP7B114U8a6
UKKpA9/OUJRBzCjUlqB9SJwYHS3OZlcAHAHMQwbuzt2Al4LKxdIpgYALbWVnZStk
9evjsyTqPNFG+19k40jVAzILXoOSSWenDFsq9IP+OdaOa/jApCtvnimD6q+se4Y9
dohfl7Bh4QYwnCdlFr6qRjE4yi0eTtRTubuTuhoApx6uqHm7AVfWWjtaUID2dCKG
n/H1nbk0DUf0LWJ86oLBT0t1trg1ZYXtJYHnTnzllBwQfbq7mY4tQW7F6qoctE1J
hpqfMMW6SzUtHrGnL1z0Rc6ASa6MG9Ib8ieSbDkW473qnA/22ve2l3Bqfm9STOu8
P0J/y2lkpnlV49R/Xd8ung+5lozq49pIr375g9WmW94+SbVEQIfvklvjju4HIfBm
vy033VAuklAp4Fw+oAIPwXpRbA3HhY4Oc2POmmsN/4+4IXzlXbG6Xzjkc+KJKaFl
abXlNWfjtE0bpbsu/ZuXMmfOHbRZhP/4WlGElR+/3EM/EHFTaIqBc2bAs9jHIjKQ
ljdFHb9MITUDYbtDRe8TVLkzPopkLIk9nG/WSZaaUaSrnzDxS3qDOx/4VzRUmG4R
jABkD1Py+OJa2dx4akaV0uKCUa2K9RouLg6J021RWVcwyz0i1tGOjE/ucEp6FB7I
u//5pA2oSoZdfoEgEw2f8LbFx/pRuHpCiuRljXAguSNP3F47FIr8f95dUm9ItzYk
PwDr6SN90bU1eiilXaSynY8HwjNr4yxkxVxaKHBUVN5LBNf8araGaoh+AUcBCPlF
3aM7fDWtfup3IVjQ8l+2R5pvAM/G/2GuNPNFZ4YjE8ZKONsVu/zhFypWzZnXZbSa
wu1Y0f1PsNCsWMX9kB4uRjpwPuK6fJq2iNMdBEnkk6IXkDnEhn3eQ4NgBzeS1lHY
vf6sGz629kKF7bMn5iAgwMDnTupzl9378NcAU8lDIsW5I0c/kgwi7eJSFDABFcqd
NxKmGohT/PP4i0cLV89VjL00bR50u2U0XhE/VmEkNxMfh5x67aWk0hohXKbflq3r
l8xvE0sEs4CC1Uv6R2dJvNk63wbzCF7jvhwHx04/iEM9UGRhbM+JUKpvaIAX9g5J
c6zh0tAsQc+vnTsyT43XkjeK1AlTUAt7NHZhSNIi7LGdrIoZdVitaryKgdNgPy5A
rHCG2BzLmz/ggtvcjZZVsx/X4FmJ0lcqCM1FHLYBApCPmYWUdR57hPKKXpCAtiYt
MqTLYkBFJP3AF+WP2W//K9lgNJ52QdOfsF9zjVI+Xw6yCMhawudiDEaCX+YsPEV6
hfwQCNIUhEBly38oETHwMQ99G23LX/dIJafRiqXa5JxvunC0IMI2HcsNQ2LvSvTb
EPurdKIzpUyAFgaftuFKJiJqQKb66S7t7yqw1GlpOlSyXxQ2G//56Y2Ip39r322Q
AlAEejQ+HerBVycaFJXwiK0ymsn9ns5A48FoHzNkfDL9fjyjwaoItD0u7pb5uyBk
vrbLjMYsccSrTZio91gfkgTXrNY4q08zj5yF8NjnZrfMHRlqgNZgO+IGXc2v2CoD
hAh7a8dHZThkx5x4VST11TFkjg+6DmxCrv/tT/iU3dJ4BaRd3SgmMu/LypDkaXPM
G01FZa+joGznQE+MvoLkeABARWXCwYI2K7eV/X+9sHs24ziFU7NofVoUmZxWsW70
QIbj42uFuHUW5dyvJ2orCcUD9fYdvsmhKZh0vZMIEf6H/TRIh24lKzzgB1EjZviX
qv3jik3Fpg/oXyOyCz//BsAy6L2L+WV6BBNjV5B/WXpzs+XUh7cDWrG33U8+2s70
WajeTgaTyZJaVcLrSnnnP9O9N4Z71YCwjiecWtU19UrlW9d/7ij5KN3twIGfN4Yk
U5BvXC4Tu2rISHDUsixZ4RdjpkGgHSLYNFQIdHwP50k3+it0HSRNDJuWfwFeg2xW
1u9bIMR+1b53nCAn4t1NRtPJ0DWsln5v4xcTleugHtPJKQ7jjhF70TkIPDSIUWeM
D9LOT4v3ibzO+8NH3702cE4vgIUmdmWhAmwHLr5txV+eIXgAkUk8ahZwnMFKCplv
6dp9LUCe/xqjtcokxGLNXr6vhqux7kKSi2h/QwwPP2m+GpMS6AMlxJa7W/H0m6pK
D44ONPLQNCfbuf6TKyhSnHqqplb44ABMV+NNDfiaq8C72E3CJ4wsjj+LrfyH/ed9
T80PGE5fL4BK5cty71+0n0YKbPb4WoSodbNq8Jqi/fnqp6FWkWu30hloQHedfNo7
eTiwAim12SkjBvpdpAWM6ZAjZvDZyo6u3McQF5P6G+5aV0+fVqorlTiBRaAL9sSR
rp2QBcOJEOEaCwO7n/MXhmSMlo1DHw2xwjEKJd1jkLVIo3SpxNOtI9Lu1HoMaKNG
qz/fXZHo6/akp9BVzeBHmGNkSXbqcm7rhxKJsNRqZHi2xLJfLBYPTj0kQO9Ms2AU
I9Er5g3kKGFxVjfNRQDMaiTnHqz/HGo6mKaNkUKxKyFQlBtT19KxQLUHWav3mrTW
iYx9lyE8MqYSUA0qg8b9QiQmC1qtJQeBzatLFeyNko6k5YB0E/DB3s1Ub6c2onh3
joAvvO+fq33EfdwwEjEQzyMwJV8wc3yPA6+//PXWK+JI53Fio/GtwyGFQE+bP+3p
5j++gh7mAJxtk3t9jnUpQRyvRKNR3UkOCvsw3+H8ybsy78UB/7ipLkt8POFP6IyN
iGEQjVeNfu5rmLIHlfnDBIueBRjR9xS7yXwNPOHcLXUBYhF6g77pkq3BVbliIwM7
43WtY+c4h+qd1bVSyqTkqQfvwFX24/E/O7tazLIuNsSlYm1rodlsMCmrrsdmcuH2
jsHVF8YzIpsdr4uYD0RJOoqoImFv/jHc/dUcKMLL2Q81yB7ZR/lMygCQwN00TAv8
OLipkTo87tRalc6gkbBki0qpKbKTDYmGPScza4ZVnOlgVNnPAMEoqBZHSIaGTAIS
vrfdcdczSKakXfnznBVw3XM7FY8kGLTgdpCQLSojdWjIWXeWCJczXcR004Yx+JcY
Yp2hL++upCuYOEAMuJVHcbe0QrHpAJsSpeMS8uaLQE7ziiE0IJasraTM0JiO7qEK
RRktHHZXBAbMMuv7kAYaqRAtxw9b7DlM2YdscQxqC6FdA8CZhur++3yhnqgZzKEx
owXnZaI/5Z6AX+O7h1OjGfa8Rhnd4xfFnCLtIgy3q6OewzjTGICELs7C+QC4adD+
5c9gKDOiUC9QLcm59e/JWwdugKhinB7flB542VDg/PIIDzpR8CGg50ZA/N0YBpHa
FxOefS5dC8yO2uB8oeWDvbIeysoNW87AdH0NttOAJU/peCcu1KanAOYtPaMZEiiq
cbTNQNpn5uoxu7peHTQDgQX6AoLuOpJlRgFluUEmpF/AxP7hwOrTQmKOHCNEt+NP
gDNWVSa0bFCjEZpWLkmoBy9y4yT5pJ4JxP0p+dding19iWzfx8hXsQMj7cuKka2H
oVsJ5+HZKcaHPIRGfcJShFolok2JdLDtyKO1kdI/pe4v4eycaclkoPr+OJEq5RsK
shTM61Acit+R8Sq12Whnwh53k8zDJnd1HnMUR8esRf/6lz23LYgOJHZ2oQDTlODu
9S4hBzaHjVaOJJQ9QfjXM8STyiNQZor5fOIoZ//isbHlB7mrbE1X83G7+NnlSv2r
TT3LMLhQVCTgptxFfBWTH2rEv14Oo+U9zX47nRHS7Hnmj+rVihuHwxpASH4u6H46
d1b4wNaxu2G+H0X4jfi+Tbwp6dMvqGY3NWzj66ooQDsGsGK/YuQFDzSdlNq7cWr5
19VuPsurPF0OEFB0xsZWu0uPik4p1MRgTprrjZNuZglGTo/1lGaWdSxMJBjBGiBT
BzFhzfMp/HycC6JlDu+pyDZG1yBZ5oqQokMv/UBGv63sXc6ToUZcqiX6SYJSYivc
pWQGMdxYn/eY1WehtfSh9tPtn3KmAtJItR8xvxt/UX83gPpFzgtEWXoWzAN1dx/P
SLgnB9/zzD4+VbDiQLqXTY4JpK9NvU2rWH3iL0AkWMctuB7fLRC9hfpQKi1K5iNc
hKPTnf59sUeottnv0if71Tf5ljmVEsEXhogJ9SvmSUSG5y/parZq10FtS4ziqnAY
cj3GUWGeWFmcsLU1C4eyUqp8EgDcZAgevMBz6r2yW96UpsKPxZ+a1AjPZlFPYY6q
6Hj93M/2W0PoCl0Xz9U9zfEUYNq3PNCdoOzsq0/bNwa6XR1qF48XdL69JJN4E/UO
b0n7Ugy0FxgeKUp2oqNAcdux6jBJ8iJRXJckCXT077zMoxkZDS4PwXTUsL6eVgfe
Mf391SUgZLxVSdsOLPCArYKCtzXrZkwGWa7CcUEWPUtPOSj43t1M3Zkwq1SeRZAZ
OTHjFlmovTNY9ofKo7Q9QC0k9KQCIqMcD4wU/Fa15oxZdLr+GC1s47fiZb10rcos
lhSIfJmav3UNUd/P7zZb4IVM1rn+GLI3o+sjDLZ2+UgJ9Npv4bDYn0zQqlWXgeGn
BMCMK1aW1XNfQftikcMtJ0c8HSYgDGIEvDlfxnUZ1mdHa6cTv0pd/If6irzRBGfr
Qmdt8ydTRdljiCk+eIL4TrpLMsf3ogijJbieEiTZ4NBpVsizV5/fzeeGr8pt/50D
qC/cC2AJzfocgoflzo/fszRDOLhq72+FIoUTe4G+yDX/Mcf2LVpsps7lST7s7HuA
o3RjSsyYRoXZgpApY85KrcORpO9jWLS6e3mRhr4rzJd5pdM7h1wfNu6hhUxqMMPJ
UqJ2D0096DMFTR+PRf7klQVn/a3Igg0ai6+/Hf2C13SAgyFzSe7SoxulVJpie0Tq
/72sUafTa1/MBu7KU4yZAcl/L4qewcVW95VDi9gWO44wWGe86v8oa3aQJGJj6LfT
tuDHjxgJ4s41kzVs6/WiIGcejcp23hCHSERqqWVwSq8RxJyQPd+4kgZh2KE7Kzao
AEre8qF9SL3kHPQgQq8pAYsaA+ve+2zdYIpRwd/8HxQWvL1MXUfZmbg899RpunnV
mmhHyKdxWOFJjyobm6xWkCqjA6Kg/AOMoeDEdeWSqWD+/izY5xGI8E5grKq+dFZW
x7xdwZdJuKLCCAIxVMLBL6jHULGW3XcmlTbWOAdmGzDijRcaJjiJlqw/wUrEaq3O
X0ClbM5/lo2HfFIcgiTpAMWOVGSKnMGuvnqdAd2q0+JMfNX9xvkNdGkyIcWEmzr5
K+KDIJRg2g12pXojRoMTDGhnjZFgaFb7IX0ymdzuiuZjTt2uokWAOX1RsI/oBjqc
jLb9b0fpjhbNioV47rVEhTcRsVQw85x54S1au1Wq77ENKEhZk7w4wdshdF0MUgG+
HDJJhl26DzM0D9OyfwSFYJfoyIyXd3NzU5FohNuE/yojG6VdAn8+L/z8/MdQ3sWn
4awgewwHqjhSKkD+okPnxCYV0Xy9ycWXsc5hKYpMiUoTpqi+rF0vWIRp/F2B1U5F
J17KwdYRsm9dhdSkLBnmE4kp5Ek10JXDbzVG7o7KmQy9LrnhCRRS1JYUOpa2r9mj
x/9jd1uVfThNJdISq9jS2pb+9qu/KK6CknXmQnBfyvI6qua7jbZFgeZsI0CMjpPo
NbtpcEf7m5c8uU/70oCQohpHWPoyyncADn2prfEppdMJdEqxqSrgrAgqgPIcQiRH
QxY1XQWEvSfFck+nm6Hxaol/fJqWi0vPhGZQ1jpaGm3qF1W9HeusVXpHWUMyNrM1
CXmDyfUEp46duClukVXbhlyc3KwemTcFr+NhcaDLMsaYOSoWXzoqwrNMYXkE22Gu
4tG0ALELSorXwVqRLvPWr3Z1W67wi17hFoBJIHWVDbXO/VJb9d4hqI/xo8Ir/eS5
pVkRPXLanV2B35dOLcvrTJX75t0LWYjyDKYISJkOfW1TnQ2MOZqR1VgAk7FlPbcM
3BFFNBIGzE6UQwf6L/2CjL1hrABx4p4z/4p/eZJaDRdy4O5gK+oCC9hdW31DGgoN
0OPbcV9mLyQrDOaTjXUa6v8C9kze1e6PoLejfs0aAcn/Z8rshUEVoQPCg1uY7sbu
GjGLQ0niV3M6AV85I3+iH2/gxDySw5y4pr6gls5/nLw1/we9DK4lIfHYR8MnKmhQ
482wp4WtKhH+TMxnCBrvDPWD1Xq6qnZNeslNQK6M//g4KNJJdbgBiAdbTnzIWUHa
YbjxF+O7C0PbLRIt2Fw8c06SherJtduLuRNKb6ui4H0d3jAOEDUerkNQgubIucfn
guLmutenu4wYtDnQGiMcNeuTBkz67sxSCpJewLiUVU1iSPZ9LIbKuW3tMsJfH4be
devE5WOxZh89okUOto8nqCQ1GlF9ZJ4Z/2AB9OCbbqQUoZzomvm/Qmke7+SdU0JF
eAAQNJiMLVV8LPIFNMsKUO5PuDNU7RbsM9d+kn8p5lup6Y4YqG/wiElnOTqcn3WX
z9L7U6AAdTd/qmRQidP23acwQ8sVPLlOaJS/5twQDBo8Z2R2FHBoyjcbSRtz/3w3
No3lMtruPvyucaTazhLgf+Qq8rEkGQZnUz5MDo62mXTvnOljYTaNG0WlMgsQj4mR
n9mApb9R7mEUVt/XmDCoxgu7ixQBsj5Cl7OxkQ4vRBzj297mOcEShgJZKmDuM3lk
eMOF1z262c3+BboTRAzIURw8dPp6fREkL2DdngJD3uu9yOAD5fHIoinfIOE+Jx6B
G+L6TNfiM2xyfTz6M77qkY7Q5CVmTswCIR3TUaOj+PNuD10V1+4BV1egCECVgku5
`pragma protect end_protected

`endif // `ifndef _VF_AXI_CFG_SV_


