//----------------------------------------------------------------------
/**
 * @file vf_axi_slv_hndlr.sv
 * @brief Defines VF AXI slave interface handler class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_SLV_HNDLR_SV_
`define _VF_AXI_SLV_HNDLR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
E1AVJkSTnr1G46RRIOzVwomSaS2w0wKuFT6MPLiugIxweSyWKf7Lam1GeGHFUWsK
PaupwTEragDiVO6k46YyAT3WfnbfKNV4pC7n3zRtP9u03avhcJYvWc/bxrKP6/b3
vp5UN7tR8S16TPaE/Z/oL3x+j1P2b+PU4zN00U7s/s9bom4gqus0JRU6Vi5MQbM0
yw/59n/pu/e3NLd8bkUdau2xiiOn1mMFD5Wlf0kKfvYD+txwddf/GruABr9V7dD3
YGEVUGdmGUjRmrFLsVW2D5xI12WUrXPQvVQslJ2ZkKzH9i8VRQWm4U5D4/2ODui1
opgSqM6dZ8NCnel919/sYw==
`pragma protect data_block
3N6ScbKb4TLewrtl97fVRQ+xHwxGPkYLBewGsOyu2jRj8rBpAbVKfuJwSyAIEl8k
Xsc8OFf8DFdFAE25W90qktl9S7V2NDQ818jIWq7M7Y16PMNuUH6tEX3sAfXnuN06
FJjJZqbGIwtmLry241rnQJwHdGuKYc9SiALyUOrEWIyn0UqB1641uRgDnWz4OLxk
vKJvUhImrjFTlyC8L58/7pFE2kUXDOYnRU62M6f+tfg2UXywfH4QDQ7n3tf3rcrO
xV7fAxiJGpn4II/bCTU2CccnzYnCopnD41gpkOBqs/OsDTkykSDR3/xvfgss1SDz
A4PC3yvzWxpJdSIHPN33Kvz+BWyGjTdWboSpnE+VFihvAQqfETEWZxJb0b21ZNLb
IhMXPf1rjx9cJp7+OkVh27wbmgGoMaIs9qBNkSWNR4OL6pXCq2ah+9ieNa1iCAcR
nqh35WvLknMifO3MWqO7uqsWICZErLag1YR0N5zxetiNDulcxosRDw1e+8NzCulp
KLdk8dVDOSlDHaNIqLYcaQQoV4t0LiAftQlp5cxxIrpFnQwCHzeb4ZFZ1J4wJeJx
to2EpwtWY+VTkxu/QZwJXlnJfSlswFkNKnnQ20A/dMjgeZ61SSqBCUD7SzjkUELg
uP1Avwl7swMNfYF+8oapUUc89qObLM5CAfr82mAoFFX+poktkWoIA6wHcrv5X28w
AoXZw4y7Q/CsbFbupxSGMoLhUFgdwCq5+kWAONM19mo5nkm2Li3PIS/Qk5r0Qvdn
STetM5SyASD7/zlGCFjPh9E2KoqRJFLtiTrZ5B+tdClbzCwSgzVTL1L8YQl5jPRM
Urc7Ww18YOfh3WQIhn1mgq3qTJvkc8yzpTjzabAc5VHdEW/Ty4RPamffwXTIFgGM
qXB7VIGV2MtX0JapaWpAdikAdRJl7qmgMaKjrRnINeiezgREW6Hq+EtZv2hKZtfB
0WRl8Z6I//T3Pvrg2ACBXya77286EKrSF3lj+yztMB3oWZTGoBUhx3icSOhLNJnN
Dnzct/vTYhEWkZlXHEHKa94U3F3pAkgNJyjkrevBWtUSIaa0TR0Y6wvYNVMLF2Dj
WcZxLtI7Z15GaUVFtP7XmLo8clFzUpCuahYy7ctEsHqk7i7ghrwHlsxIepWJdBNw
Xaw14XZTFh4tF6sse0ELSWYNQPIyejTdM2jvd5G8uTy3hawQ7eBWC86QIo9GQkD6
BzBWNdZxca8Zk15XnH3VRy1cOWtxErusGkuf8nAJPYJPyHmt8hz3PDyQ3nbgq8JA
vO5EvwedDLfAv6yvkFkL6NBPDhxL1CIEv2e8qwXKIlfIpn+IAW/TAA7ld6acFOhc
92fPReYpvZW3cL8hpYDi35sfYJOOchhErYFt+8gQGDV/UWn9wqqMcrttzPLyr6K0
HuVf4B/9feKppXoS3mUCt/7SnFIj30MUYXtWaOctdgm8jWu6RblgwXhNQXP7Scmg
UbPLJdBOXjVHT+iMrCz++eRJNlowbqH9Ece6MnOIzXC1Lbzj0DTvJXtisIuWRxb3
acKN3I0WmzIDTybg6TWzbqJsvQoiuJ2nIhNArRiNVJ8RYgnm58hkixoRti7u/MdZ
X8RRAHsR2ej6xsI8H34ZpE1A44s7G9rDl26h/rgs7UveKdTyNNGV8cdCMR5WLY4L
auoKn4dlBaQlbgfMsHiwbhpZpnDP7fGsToIbvEm7J0vtTzVAZr/XTMjVELDiKVhP
dxc0EOdNqqhYJx1ZmpZG8TVAVFHuMQuZdddtlYy7eNqnQgWWX1CiGUsGhUfYwcjI
pzOZyC1XBcz0b+wq2cwJeRpsfUo64V4tsinxw29039yIREhQitWi7Azgex61UKkD
pezeap3SUFAKk3EeUn0N/vzd0s66NE9Hcg6ZB80l7Wk+q2F4DUUmG/0MhNmBN8ty
G5hVyEz93En30Q6c1uu5mLoMPgyZZzc3Kl4wqZ7NVRadGlBv3q3uB3UQ1HlSQza3
bRfLoLz5Wb4n/kQiVdrRVBIZXhBH2wH3O4iBpNNCcpiKWRVh7pvHW4AjwrprazfC
X86T4zxr9ujcQRVTPOxUj1wP73B2ILqbcVr9WauoXnWjpM4XOK2TtTg0bZ10LwCZ
WlT9ekHgA9zMRV8+2hEU8il314SIp/IvOdPZZGtvKYf5hRPzX9UrIgG+9WHNQlKW
5aXw9WotVQ3hhKgmirenZhX5wB9BkB6gPLTJv5j35lvq6vyRxugHIx+qc3iRXN1I
p4KwEzgDFeHniLNTIpptW2cUqwzi5A1iNdo76dSxVW5EGb76waiLl3QxVYMrDjBH
A0SOkGckmPjEQv853v4uxRyGmFCpEDiPyvk1XScckf7JLLKUtvy/oqIHSJkVryTC
EZpanqdLUrBeI5ikC57NyZF1KI3iuiEY85j5ZT/GjsDZf2pfxA0ieX5tKnsy714l
DMC+NiCmLkNztIRSezvGyF/nV3nAGk4X5v/bfh8GmNzk48UoYeDecsWnHRt2jG1A
h1zwa8gynFcf1+cxym9OM8SJq1BG1EDicHClWj+W4c1p5c8v4PJqQJZpacOO2H4a
7YfhEo0oQZ7dS6W/Oe3DfKdYnwwhFEXo44bDUlw8dbCQgqnIWsJledtqSfrc1PxV
JcN8ktU1BwTlenfj6w5+D/UXvAvN105CXjKJdXoMC+2tCJnOnT+JcF2NQgZ0CZC+
716Y49jE6220LIIYZ9m0ZWq3Adq/0Hyxo4l2hU1UtsNKzjaU19RjHtGIOuNIbk2O
GD07Er2OplVQ6TeL2R7GSWZir3qUW23yM3KuDECg2SBxn6pdokIHSpTXc8fSmTeE
ejIkVojsbta/CqajPbJlRKZ1hQRgqXW8DJohO9SUDo35tErRPjeSVRmhHzisxIVM
pAsQkMXKXIAaYqV6Jl9o3Jsw6n+VLag2VXoNv/vltihty7vHWoVsNz8EkXOBnpbW
rlGKnyGN63QB4LX6wMSREttXmaGMhphoKlFFhtTcWDtluzujUPloPabApUr5fzeR
jnUNBP04kt4LVfmPFOnPzmRXleFGt2ov2mTnaqvf5OGmiOlKcThp/3Vf7y/mWEKE
vPK/8cYoPq/vL1vV0xfGjwuVBXy+fPDHEGS3Xf8LYi0Phn2CwoovBFbJTeXAaxS7
SWlW+41Ad1tfZIMIDbcFbcq+EaECMn7xq2okBLFKu1Zt2kOF//PzhmADFSOWQkLM
fdkLgInD4kwG6kaqS+iWxJ1va+X5yQmTw/sAzBC6n17tbWGyM+89pfVAkilA3/CY
FKRJjo/ye8FLfLZN7kylwaBpy0diu+wcWT2cWFmqYEOhnGNUtsZYDgVjB10WZEUV
GX9UnxkPagqjGeqoDwtCpUaMh/wTPUnH6P6FH65ya3rad8eoUFnwcVphL0Iwux1n
uhZLJFcL1IidDkvLHzyzxNDYS+LTE1i6MgQr5ldeLND6oJ6YY0qpeQiYyQqpk++Y
F6mDHBsC5Z3TWkNPe7brD0exUC5Q3FaxiUaTeuBMYUmCXscoI2320P45H3iTdnnX
EHVC+jkru28C3MwZFPBrHGG4/ueGC1FpcUh112linKz8ikfhRayaJynghXISd5DZ
zdz1DBt1/kwqJWPlKGbW4LIO4FouPhmzuxbPo2S2ghEMNRBEVKUAmC+x3CExfmt3
qnFF1L7uET7+wK5vy+3zWlyvKrLufXZsMENNwpyleVt81ifZFivANhX6lRbJOI9v
M7KPbZwJC23jFyhkfKjILdd5IhYkpogCANWvcjWrq+GGTKAaph1yoUXb9+X7Ykse
AVLQAoaPpw9mlglCnNj/N9ItA2cMoNcOz1ODvwO2I4Ynv/TkDLJxIOS8zH9dCGR0
ZmJTd7+Rd/sToANUGA/j2ufp1Q6B4SqYXc2BemjNygVteNHQR2KdJrZwXXe2IANS
Jw2hukZsZTrBKUjnYCBXnElqzCFCKg/5FEnHBmQzbD4fTvdbhCyqM9xKl2OXM0XR
fAhV0JuyzINuuB488WS0Sih3at/7UznOrTqpU3jsTvOKVEDTDd1FxNqE6kTaSNRI
nASGzVqhDMkHlJ/dLgkDJS38058DyV9o8Uw/bI8u2uIy4+rnOn2iVrYIyZmRzKsq
W8dMhjwvGShHotM4TUf7X7ImeiOY508v+HkERUm+L1V3aJabMPOocZgrUtV/t76f
Somwgab+tHppgfUNO5yqbDhfOHaRQURGBB9r1VzAoCxfjmide++1kHoMV0dkawf+
qnMEcfLM8bFyXB9eqvz+DojS2UlxncVsowsYpriUVYDSYdiPgr8pcUJ4WLQkirXF
LCafZ7R3lHbwUUdkl/y8F40aIiOUHJ8hclzhP8wTPGkfQM4afYm/KOLicnHWWZ87
sXLKmDJyz1WJJfjCrAlDDlOGtyBiOXwRsdb1+NB4QGHUTe2lY8i/LEutu8Ob1aBe
dRb2A6P8HjkACMJMczyHKLLAAZFYeexa1s9b3CWUnPQ3uuHDqDXtyCCfzbvgt4Xe
DCKPQP5U3DY/O2U3uxP+LXUnr6yN0SqUf/0cs9Z/jwm6LhKJLeNpU+gSRSOyhmBM
j9m8U7smC+Pj02npFyKHcspCOi39jeFOKITe4J1Y4VY6m3e4wP/XaJ5+cmMH0cKO
EWzW1A9D0HnMlBPLl9Bu2OgO0AiKnjJAmUZcTIhyu6Q7feZFS9qOr1MuXt3m//1Z
EROFhf7Au+yGmBb7YHLXV/snr2MoDdpJzbQuS7TYHTWWpJIaXFGJO94cbTWWOJYL
IvbEoCU+Qh7LGHs0RxE/TR1LDD/bIqB0CXvUrSA6Ety2zkrbeOascS1vkll9JGkH
J6bNJfwyx62SFpQUTy7Y8qSheXl5qVD1wJi56Y3DQahX+MJSKeRqf2UB0r8PJCyV
9t1UXvpKR0IiJnU9SRDkTPDK0cfl28i9xAEElBa3YESkm9z38piI+OYIgTKkSI6F
yRq3EHnH9KEO6xBK/senOVnk4gXrd4EG8Jhd3CCKxCJEvRJ+5MtrbaXU1e2oGPY7
rlG/n7eyEmvPj2lGndEHTrRXKsxlgwiuxXqPSg5BR/tVuSNMQqcqEIM4++btdM+F
mC7T6e+J4mbXVhdMtFldtE0s811lmNQhFzVlS3+oU2vEMm3T+8IPEhiTbMr2EMDI
22CznGvsn0kq6TTBpJs/cWkZF+tkbIWUA9pZT55gfbWv43QLFaNzOChnQpQ5flKW
6f5NBbJ/ikwkSJmwCUV76YECbahbv6qgeQwZ9+2HS/TFPAQyLnf3KE5xVW+Go4kW
wPrmIzUYX/ujzxki0/gVm+YlUEzSj/hqarCARu1yqZw7b0YRseyqamxJrdBngKup
fIoGMPd518azm4tvDmt0B6ppSOq7AQEzVcpCayJnQRZQvuenZKirrjiEF2QtuUKu
IcHllRMBYx3RO8iBRaF85yOM8+T5AXOmq8yIfeIsAMatQmZks3fIUvn7Uqbm5I5V
WMDa4aNcSO3eQmxXM4vhfqLD/aqRYA92LT1Wlj80Rp5dq34CqUnX6qV/fpwwCJXO
wAqTStlb+ztmOWVSDcS9ENjnQTF7f/eiTa6Cf05aGXbQRqb+g6qIsbSik1vsoxS8
nya/N08oM6TzAbGnTxb8sEYoFBuJXTNGZSGqPcvJX4TlIVSsubNeBRRDNzUFE9F/
N3LjO9omVA7ImpT0Nmyr9SxhM+aKI03vvrC+GOLYIOlxVfGseN3QuHvCmxuUczmH
vu8BhNBdVRYWxRg4fX3gsDyZ1bgUi009VZtvmtgk3UucSVLVLQ0geagJDN/FlHtl
vNqFl7CIPCug2hiYOaoxMpEy0kOxgFXRu2WwMfXp38yRiNUQ9EJdtnUL5ObXCUiQ
347y2qrxKUCQMrQlN/69NJm2PNk493K9xNDvhGHm2sumRkGQW4jieaNhlKPivPvX
15+tkqIDopoYeqQwX4gfmxA3v28n5Rm7FrmLkFxPfQhE4s2+KSgfFa15aDYHv/ag
r6slkWmcAwzMdaIRgAKmu9gZIE8QiN6Q/BWaYG+x6PrC+5EsIjiT1I11j1dgcLkQ
hYaF/EPp+tC854pO9F+oVR+gsfKeM0UlD5jVf9+SqF029svzaVW+QikgkLQv9ugB
4QTUOue6T+44ohYg8MQ24ZJGa8IgW3ocnNV9gyWtBC3nBHMrFOjB/tQF2wOB7OIS
98xxKyjcxuPneXazkO5jnChlsNH8ha10SYkwvoLECDDEiq88cA3Bk94bXbDBnQBt
k0BSMMQ4ulNwHZ6UQSp8gzq+QwbeUEsKQLP+RHInK+rifw3Ir9IJXlXuXqyV1C8c
dKQp9wYm0I8aKGDh5Rr/1LFjTkcdGXhwIeRUl5S5WAfIzgGLBOsAL5pIDK89eDVi
zXnelNoV5hKonYmvqKa90tyDvLKjC5B2G3CGazFL31IwYa2iqHGbEeNAIhv9H/88
BQuZXP2CnCG9Fyjelu0ZR4KU7Uw+7aM1c3buAn7VWwkGTUwQzuqsZsjBfzglfH3N
AF1nAK8M5AjC6iNs5mu4W+Bv1AjsBmhV4hDjEtgDgKCMx3xogM4pGMxf3oafCzub
mCeUo8t5Kkkcz6g7Rm5SS5Pzk23SIjE19qXgVAmFqNyAovSc8EhcW53s1kEwcZwN
97tjxErPA6JoJAgKTpLXmj7We2mk/pEOdu7cgTtZ0gXdtMhki7P7BG+BvKOyXr1o
pxecfA2pcQKVPN6pCWraeu48hVzTdRQd2mMfc30tfb9QO4baoJF2vKefEa+DvNRq
9vGkCXwT9Qaky1zTfD9Wsk+2DZIvjtyyduN5ISNtJCuepsaTCuuclmW6Sz1fysVp
i+tabYczqtmYGzlxwiOBVpfRbqBoe4z5LqCvsYUERNkFzYxcy5oMcYTrKbfkROWZ
OgCZb7MDVqyial59R/rC34UDFcrkzT4wzCkAL95MTM1SxJlBUUVlQl6uof/vA+SL
RPVUSnJ8iFUTXPx2Ys0CEFBMB8Dx9c8pqC7n3S5YOU7yxAjgb0afeQiSettVjbpQ
SB8drjrTNrU1ZZ8LSrBA7cNh/76hJ/BgGKXYJCsmHIvvA8iV2IiL2TnLoTZiRzv/
zR/qsPYFPL8N5/jxRBdATO0vp7uvNHTkgToHCTH0LWTU4KpedhxotEAyHM3wV2Ss
BDcdoDxVG0R/B+pBDhFENakQJUI88vkRjG6cMr7uDgq3uMlAFHUvBvfUm3uiVwcq
XnPLvix3QPUUFOf8Abxehuut0qDkzy2fZf2NtZ1CA7f7XWBup9mrM+3vcng6XF+k
cefOCCfckzJX1tz9/Ll0ViFDZ3kbmJ24hFdskPoVX4OplVUQlPB4XOmDAgI1kmoq
W6tLkiUQj7anntjr4jyIdfSLUxi2UuEaviE55x3WtGtDuvO9zGo/Yf3/yK0Z0dNX
l4dBzz8XLfoiRVznhoAEeQp3JP9F044QqQOpWuwDQW3zaHhxz9wNui1Ew4OnnuUf
U2m89I72htgBTZclLmbHKJYmw/zZ339/GGq27iX3T3MR0jgsqW4jQlNWdxGIBgtD
58lfUmgrQn4o9ddnU7vphPjnVmcen0154MMOqbFVveRDuqwH5D16dlYTqmAibN+/
2BA196JGiEFc22PVqZufPCLGVc1h8VEGCZHQb8Tvge1Qz4HJQJkt/3EAY99n6tzx
1s0IichYrWURsfKKmCnpIhtZSz5E+4S1dDdOaM9LWm/yikBDiYgFz/+190ahCGpY
0hV9TykigMEJIXySq6mzzC7o2vfovGFaBuymzyGnYnI5cX6ina5LpVRuSFBRxPpo
Max3+Bxu1/aXB8Ckddb330n0Jnot1amzRGtFKQqwRyBrvfrAodgBTKdATeLK2LGP
Nd/kJ+rS3ZIwXkVrzInrZSAAXt3Bpt7EBQnLdlI68wBdb34w0AQlMApc7B6f/9Ys
d2nCt8VsMrI/q9mEb1NoIJBXrR12olVOFB4ThHhSMbEJFWi37pCXe8OOJEVN9/4d
aIV52xRnmNDLU5UHYcpBRikTaIARjZu6DaSz1treHQSkzB29eEC5K1aP/OY/u0zI
yCVWYNpgH0OSlI/nPFLoTn7UtD8o7vH/7f+L1LJmqTZEm3pgKQYG1zm9cJJv/Lza
bkbjMBpa3vBjWClMyCyrOOa8COXMAI7pgKvdZoI/E++CdMJq6kv6wPjalKGjCUXF
QKFo6pqjnEKk6hgguGlhkgoQ2xGmf1pH/ormPwddELJ/GZzMpcnwbRRAXDg0iRXr
1q5U7DW9JS9l2UDmereY4k5JxcDiU2UdYnDYH4fXCmzX6sKdSFJraKy33Rw2BZAN
PL0xNJZSO6NLo+PSJj4XkYmrpC55IlWNHWD85lPfkMEj7aiRNJeL7g1pDUBHvTD0
Fu6OI9wgfo7cu5RYIVcPjlunL3l67tleos5IJpSV7lQAGNL55N2ZTC6ZV7bNqQwn
Nexla0Ndc8vaJBPz5x/vnpVfWpPZFxn45Mybu50/yfF1Q3aaQsgKIak42wRR2uVn
Z5E9e3CGgznSKBiC/w5hUSffAyWl3iAA398k3HbfVBk+4+DrY1R07uoitTAfyKAC
j7vjqw8/rESXSKFVNH0FQrO1AythFo1r8itdkLfWRGxsczIqNu8v2eVWLJoWwXcU
6GPmBQTnswuroomy4HVCwXED/h/9Bkx0TIdxLz/bi64qq2/nyahcPuwgO0GBHo7E
6UHbAzLmbwwHRWQXvAhbBoc3S7Hh+kOv+sGSip/Nwx/1h95O1XWdO0T0QyUEyo/F
WHuMF/xkEmEJPSP9UXSfqhkWq0MhLpL7fDkMLqC9MWJtNqiuYXFwwSbvVG2fHu4j
/gutF7+8fomfVuy1KYBSfhCmx7sg94V1/xLNddYpQH9tV+gINWcDW0axrp8/Qrgw
jzTT7LOvrZFazU7Yndrn13/1ORGe9UYjs0i/uNY+6mIkl2MTvCB9xn+r7QtXgCWT
EsE9oECoJoHLQBgv0lnR4UBT92EuTU0HG7zqNOpjmddVqUXQbHwRKAVqv4O3CO4b
tY+3Um+d8xsr1mi9f55FMtPlAGGRK3BIA0gM5gz6zbLi13MZSAUbySX40P1Db1ct
hsXxOdy7fB8BSGSHXc9fE+5H4m7rv5qLm5mL5Ivv5dkaJfodrIeroAAGL6Ke7oLW
Dz2X/tUaD+LFexenzc1ONJSMXHAAlaZrujJo4fvRxOMyakqp8djpOCWwzihLJ+Z2
Ch/5Gqe3B9qVjLLDxweVyTOYckrvVtT033J6mIZtcYaPbgtOUdwiDAWw9m7wqDY5
H76X7rFO5xB4jWs0uIqtXb6wF++ZrLjmQ+NirQpFC0UrZiXjUn9FltWeDaJGX+jy
1+T4HPlkUcpQPFirMHYDda2dvogCrNrLssyM8vtIvB/Thw3UBgODUM3UeiBHtfH+
lnYuCAcY1iXvxTW92p6LK16hjUvJEHwcI9w5kcCoy5mLhbZoftO2/EucOCMZib3c
QTClikojmSq5eOgRJrY+5Lc8HdXf7qdhWCUlaABGXa8ZCgV7+p1Y5E5QwHvI9Uox
YFRcDxSdp4S1kudG2Q0NRDJ77+8X5IxfrtIxO7nvOFO+mQFSFoYTJ5U4pqAgwfDk
0jueYd5gsc1kaPLypocFhKTzkoPvL3xDVsBOztPFnZoU/IaeiKC5IhU5fnDs5bW9
vwC3q3mR7g6X+cI46UrtKVjr+LXaIosoD56TepBR+u2AUYF45WbMXiHvfUMnq8aY
tuObnd/FdoXMX6tKdA4NqMzI3uZfE19XZF7XvV2lQKEkIyMZcnwyKbWE9e9L4+TD
Sb+4pYEyAWFq/UKOFvbvFsfE9TXzTJaCTIR8C2Z+4kdD0GaYAyBctW/zLBUlSrA/
J9gYaG/ZSANHFkwCoRIXceMkFfzbCh95JAajAwpzFGeWLPvpDLRkC0lyR0g7IIj/
weZ2WwUGKLU2z7LntKTafBLvWQ7hOpFj3mxPo2aSBPrgBkXdI+rW8a2O507Qc8Vb
qoEdXYXz6hUEKX1x4PoLAY1KB/pkFUVeWU4PW1ULYnayDMc5Ymy/UGJ8aBWtQT+F
hoY/mfxxYKhuOVqMImnkyr26vI6tsLjqKmVMRyJOy96pg6uDQLldiluTAT+/1eax
1HGhzHe4LcUEu01BXImmZ/2dq+TBFLx34ETnc4BzBfGrbDkA7Nw/EDnrRBCHdHAA
enieacjGKM8qbkmJ5Q18hPCo3/aBH/I6NRaDhs1aBzwwBvoYmVxWgwMC3oK+RYN+
ZRZLFplWRtA3h+cBsF6pepK6h1zqbvQNTmhN98R22gUSpIZD1pBhiVimCMlnSc8E
ailn35AyTA9GTLz32T2vkVfRIE6MboxrxiXNIAaiXwNFlf/gyEiKG6DCW5Xu4Ln/
V4Eq/4oDtHqWtcYUYGJxZLPPdAWTyWcCz6/NLIHifzWa7T/J3ErDmnyFekmIGwmr
llN+ZhoCNKxbmnWtwX0A6wjKEREFKwe8VCjizLudZoVlGEAIPsIiRMC2uYh+0SrY
GL8cPqDYjrBJ1H99YbCz9e9VCPzPuixoJUHLLaitpMGWkHx/sKjxIxichlZUIerc
sEj4sXPUtw2ngj8ruxjNe11qJc7e3SxqOtsthYKP8jSuhqTbHJzSb0ZbNy1VVXZx
5vU7JjlXmMtMiMs13shQzbd/9YSE183TqzcyoKUHayvSxyEI8I5WWLWPDuwOtbsk
UAef+WfzVTRqyXoTlpxZoRpUm+0M0nBO7imUEpNvWf5F22Q0D2uw36E6r8w9j/0l
2thRNcK83p1uxOQUzUK7A5lACJYmbqF2y1Y0CIliiTdUafkx5UjYl2A2XJydv6AO
rwRHTue0+H6lYysC9wCR/BiQN7iX9uu2oJ+Oi8lbse5FlVseQ8+KXuKZjRJpnY8L
MoDQzFO74UE5zlJIc/YPnuhNCQ6XQCDdkwwVRdJQjME2KDhPb2zeZ/JjEvdtrgCv
TljxTR3xp4ByMPPC6/BzadAli/HiF/L2XOUUmyC/GGsJLRI4axZflMMwtG5qxMdQ
jQbb79jqI/Wo/Yi9YDcwmq6vG/MkZtpP5rW7it6pJDeUo6J/KSpZ8l62M7epp8Dn
PLWeNjOI+S2wwgzoWiBgK9hTfnZK2YHckjGib5lJx8/XE/aAs2A4UEs2uGZZQCBx
SvFVi4DFq7yBc7BE09fifoaoQfxxxAIYkQa191+5vhavHufgAnMDprTf4S2OffFJ
nnYaZsbgNBpwCNOdIoyUP7v9vvthz9lrMFlxC+0WCR7GhIsUz1y6qr751aVKH0YA
O9OlxwrrccNqPCS6FqUqCdgxJalYTpP3AzIg0WbBuk3oPpnvKidShNCkVxOArvf6
qdNtdZmFh7FoLW/mQ99YJwRdj5ZkvE1w60CoJfjznt8iOf3idrM1BrLMJ/SQVM2d
09H/ZX5fLFgL1urt1dtMpRElfCA4AL/Q+JUriHhmo5tUeVJO/D/S42aB+KrAyoy3
riZVQSe5yMthGSr7Vw2iq30IRi1ox8j6bTSAgmsvptUcZohAAU7YHGP1KAPmApUz
GcH/Kka/BUr10aTcp35fjWnF9KanJk81V/sfZbE16fdIntmxBniKfCbfocj1CTqv
ktx+VrCOoyi7OXJ8B76S02lEez5am2GOkEUijOmnieIFlQgRBczQ/Ih16X0F3Tl/
4gBE+dKvqQY+526rPenY2/jN66LicqOvoxMv0mTF4HDNuJQrnvOC5rOVT8W1qN4D
He6h1SW/WOr2s9XjZuvZPl3j/HYWw3ALAM4bowKbIC2asML/7N7+4mOSR1v5qaF+
HTw9+0JmDm69r/eAUcGLDy+Z9nuLoP81Q9x52nMMBDXfCvd1uThQyQ+dLco7kuBq
+JbyHRYx168ofDdaH1pO4zyaditGrxvwPHFpVqmWlB9DtvlTdHyuLjQLE3WqPUzK
Mxdm8lJr6Tz+i6k1yRxxnWszA8rpOhpJzexibsPLH0rmW3mSAXcRx6VQYmFzTvKD
wRAmSXUdaMoi5a82XsTSCmJbcfuIWiH95GxPNQ4rFzal+l6capeL1JR5O0pWmOCa
FX4eI8K2ShqfZZJWQI3xeUwHVhfeBVSIfaKiWCIdVnNGBndvcS4l6Zo6xSEbb8Kb
h57dLy7wsgpCBawCHc0EVsuzhU7NaGsz+FAzYGMpqb9tg8dD/TCOom+3/omh/t63
5lBSWkKG/We1Ht05z4ZFbuvCfid2spSgnZ4wh4kP9Mx2WqzCz3IOTq9bS2vO9RWZ
NZ5r3LPYXOgdV81x+b8fUrbdzy7tqspwtguda64aivLA11NJBRGpV/wtTgUf+in7
qyA1sxF7bct3Ixmv8SpOtMHrjmTwCz+UKVQYV2cnum2tCwyIwOt40MsmFsBPHqXP
C7zjFRHXesUCNvvLog1V8IaqUXAP/eh/rV0WnSr5gLzrjWJqAksqfUx/y8OWOgRS
o/mb2EDEmQz3H0i0oSCOvuE3ro9hM3RoukdzQ7pud3Bp7S1c4TMbu3OQl0a/e1n3
zN8t5VatVQIKwonsA66+MH4qzfSSJC0PQcoGlLiChMkl00+/9THPkvW08DlQPuSW
oqVUf/iuv4eblUdD/jzOtOEE3qR9+R8w8LqnwQ8FqVN9jOgKv2YAiKpVn97vsy3x
A77IVKeY2WaX//qFHAAHhTNi37Gk1C4enDTHVsJ/RE1lQlf3ktGgq8Z86FbEl6Og
eEAk8gmiwXTwA1vKdQJ59PU1tpwSNWMBTu6Wlbod9AKce6Grzq9Yt5y+BDVsbuSA
uP7lrEMWUZBmk+BgEo5QnkQmtDKzFh2LpNl6XjQR+rJKjO02kzwmbVszy/m75Ttl
kaBKZ9wN5w8FHjI+MQJmkMfq9xGAU1Mtc5L98sQYvBHEVJmpzmNqWVqHf5KG/AzH
L+OrIaKFWXnQ5QTvnFN3eCqgiKXIZ9uwxfjVZ/AvPgLDKhxE/e2VNZXybvBsiTnJ
dBwst9jfEVl/o6k1HzeHzgf2EkX3AvDbYlRX5yZni9ZM1VYiSdfs2eUUZbEtdip7
aTRmThvdIUpruecMd95r5j6Udu82bWYAV+HI68gJKQGZxIcuNhrIZWaFFKZg/Fvw
FGuU305M41A6ogdta+/yQREH20XaU70gS8CijsqioTPP13AXtzOwfNYZj7tY9J/7
m4UHmzg+CknT1zgnK/p+qPYuotiRyLA1CjEo+yk2PHnMPeIYwdzfaGgb465SKlZb
Qr2EMbBjfUq9ckfJYlHIkwPVhAobyZKsuR6uqEiaJJhDKtPZQLJGq+YVfk3HNZdw
AF3f0fABWil8cv8kkcIX3eDiHBYLYnM7aiVXfwXfmZB0Enptb5fIuDlqCXxE7g0v
JHrtTWzHr0MLHnJGsdZwLkkvCHHVKLCjD/qKX7wk0jkBhGsFNLyhjk/hw1PNIhMD
6uQt5hifNPHgZGGt7qWdx/7AwQxgHFCFkQFSZ0xEKUysfYdD3FJIujC1fpBH8o9O
v1KpjMXJ8h648OomDGtrp2ctFxuQ6kZhMv6wB9LvBtTC5Gjb6BRxEK5KSKwCFzeQ
ZbaAK7lbapJuTa1SbM/5KqrO7iu+aM8obhBbhB+JNFL1zx7jnwC0yyFe1EHuv3um
C5e4gAr6+ALVPEdJtGF6uFy+e7RTlLw5clZxG+wf/t3eCku8ngxWhjKU02iLmm7H
UJiKbM06IJx+S2KirZpGusAvWL3aBIxM8xUUtSR8phU6O8FY9GtYwuNpcci3BQ0t
GECjVaTzt7JjlRyAGAhy7pBv5yo6X0b9zD5D4ACg5xs+ZTZYH8lkf0KHTEknCzTh
uePK6dSoy+jqxy76KXFt56nIM40vp3CPAgul/jiaSJXLjyMXLX7fWOpL0UvmxJZb
zEFcbD/CQLXo5Za24ZsiojpypoFrBz4iungtIEKhG66s7g/F3il66GoaC1hz4iyz
XSucAfYk+36FR2FWROTnRjlKktgdaCVT96L29BfsMzmqLVuxxzdR0zpB9uqMHDJN
5o0BRPy4Dmix08BsgAo0RKQJR861KvU5yv/tTcOydp0TZg2c9vLnVLaj2/anQXLz
euKDCeiOJRSwZX4KEzVMRGOpwCWWRbef/nF34gDOmbXDUSwPXbs1MdRPppi0bIFx
opqYEkw2MFhjGa0u2tPpaChDcWC57A3NWgxeMo4bj4no+E+Q8VpRgHozFBCMwYlh
wMZVFA2yWdDOVRd51MelYuEC2lAybrz9I6pPi8m5jW90fY9AxmypxnzM3xLAU4V4
iNn1Z39t36hv7EE9YBSwgDqDUnDM3/YaVJOZhoyKAPzvcW3yfH8AKZW+awFNx3Hs
QqOXTCbWLbQEFnuu/kTY/EGNZr0qzCykQKUI0wLh+mUEP2dcSCPHPOf2CkElEJAw
2xAqiSxoLHJROyxE2PnCGy5gcX/up+iKNW4WxlIYAAKn8/kDYFoeJNwKryIEoR1q
TWLLkIzBQLHMvy8bSB/XuqpGm2B932Hq6/sLEZwd257P9ci8VTS7MSRyvAZDJ5OB
sZzairgN2AJUsz3RHUCSeYr9dBriAmR5yMK9StVA4UQejcAbg0X6HVxKPQYAjsnt
yY2ixag/E90Lh8xmHuXghW+4tM+E35kK3vBRzAM3lws0kfoCWQO1oYIkPzVNafiK
3+PKnFiZnKPdq2vPI0HSTiDngRSiX8gQPbS062LB3c9IJJDhbiJubc8mCmCDsqtM
QxJpOVMNYjeeWvuYEP9WeRKrltTbAiwpeKRlkGnVtqoNZ+E3AeqmvqmA4Bd6ZlcD
wRNzSXS3FRyoQ7lQi1hynBYA+g9+FTU5iAYaMP4jD+wSbmow9iA1RMioKWFLBhuZ
Q2LGM+8j2RAD0JoEmJ/qlUe6idgpV7YdPSEW5Yek03ON0vgmIqtB2bK84HLU/Dyb
kwvN/l4vV3fm/K/lpqYk0z0c3MLbwtyGSnV77IXz+zi5DpGytBT88tx+GlI6Vws9
tLXnNwjjgjbMQsOu660Px77Lq7sMTA/W+tXS+6N4eNEvHfhj8xm50W5Xkd0rluuP
vQowNIpFCNXpJUZ43j8Qjqdr3roQcIrQ5WuDRmspQpsjpksyok3Qx06/WO6FFB/G
fgcBmTbVntF8QfcRgw3Yw/Wa1pbGlU5wpFtphnsMmvteyrmBlM4rHrvbrW1GpNTD
53r4xi2rDqHwg0jWRoMgeBTsAJFlq/ct0uF23HO/M+w38+8d39uG9xMGdd0P44D2
hlIxTsr+Sknu9Gl3yyt+oTE+2Kvb+roEF5LOH3eRtCqrFtTuvGVXgmYN4IZZzAy6
5TSUfdqpNQLU1hH2EXnshKv0TaAA/2UgPJC7qmdWOmNiNV2KH2USU7pa0qBwT5xv
7CG4gJcj3k4I6Hm8YKT/+bCuv1Nz5+/YWEB2sI3vjh3vZUrbp+Rhb77c/UTaBpuW
c5FLfPTezmLoh5Asi8E8h86XJpgRnzDUp6o+J3bBICMEiT/TSRq9jgDmUMhAdv4d
3hbGpkKkQ1ryvtOXt/QLUn4bHKIQp1E659OEnwsTJnEOLc+aL37zi+ZmMZ/8tzgX
89zr/NOjLqf2rCwXKoD2hU8Dd2V2mcoZ8byIsKSMgl7yamEhEg3pe3mG2puT2+Se
qc/8Zl93E+jiQ+CbsR/gcQj5pBk0eUUv4oEx2GLgk87xYwsmQIQ0xeO0t2+rtLTk
u0FSY/P7PZz0YKC8MykJeEnxo/lqW7elDMt89VdAOo/nHgRfjHcC81hy7PPmEzIW
x3WLsn1BK49yJO78TuZRnyEadeEW4TVF436lPnSpv8a9gSRIdrjPoiAQxFRkrYtC
cuvW3DZWqN9pFj+/XEHJCHj/OO5rb7IdYd8dHTcNCnuhYIpT9eOwgAAlDKxemXVT
ERONI/JaFs3RWlCHhqBBvOII0N70yx+vjcfw7EWTigjMSBdLzMYi/y3P3rFX42Mn
WEuV9frJY4m4liF3TxIVeotxA4ThNr1sHc8ZPX5aC6ntC9ReQW3qeo2rIMrTGnVk
SFaN6HbbvqZ1p8XCQlafzoEvASWMbqJL4oLnVMTRNP2NK/6MP6R8BZfJYwOrBCvr
/+WFtiNdSRgyH7Ti/CmIvtuXiu50jUVWEC+Xws/dvzXI+jwlbzvc98b1b4nWiTGg
24rSmfj0ruI0xuogxbSarsjzF0iPdqPHpgjsrcWpTGOBI0mG2NrbRsjPIvK2L0wn
RwzAbnhGcCkGnbOqcS5LIZD+SucMBcedna0OD++m9OrPAvVpmihUuulknL8DqfSj
4ek81iNxYLaxaLtL5CojdBZ4dMxMZXbl+vNhieLmtU6FT5SRPjPTOI4R/JnwsJes
js1InbvNrIRSshLNOP0kX6nQ4tUeqTQmtL93WEa8qorPuZ8AL8SdgtJisoSXpzPL
FKOiva0LsZ2lKKIaoLHdfI5OqE0KNImh9hCsDWFBGhMYKsUMuEt0jeZQQGVpbl7h
1KyKi8htkVLCVe2ypHdKHnEuyhvJ/T8p7spzGSbCT/WkgBgGWUdVuAvlVnhQHPoY
s2i006zQ1HkYoUK8TfundTqevsrtUvhniPZZ8U9v6OuOZLh6xwXN2Ex8U2hkgUhE
uMtiApgVRhVJsuvon+JdTVMy4k/xylKkGsVtRUFUxBigVhf62BZ/MbsUA+mqA9U+
wFpB5EatwZXnsQn9ACaMmfqHy1cEveASMBAMBI/A7/TYoUxXNfPdAUboUgneJiJy
pLaJpP+Yycr/sN5E3aw+1q02mZkILT4jC4OC05CVUwqIezIXRDh4l5VeH6Ms04G9
eq3T5fHLhOHXHKNRaMn2NQdPpQKQuqfzFrp8CJ04GwPlk2axBiQmaHH3hSmM2vAq
YI3g9fHMJ34jZ3anHJJvvnRcLVy8GW9EoaWrJsc1aQZNOehQbjzE67BpYaS3cnhz
aT5I0ceS8y5yBzwLfnJz505jk/fI0tIu5xfvT+Hl4dZG4zgcTaRmTKZ6B6QZTskL
oE1aEiuFndhvs1bTw/36WACtWSiDQfqzQekqv8mPht4jkiAmARZLpgbWYHSCbb4/
Nb+npaq/i0t9kyPZSV0972eJTbJ9jHTIlNqF6D93zT+2N4UHziBv2pP9mUHnib9x
N4UAuHw6e8LrFsMx5lAXrUV/c+gQZbQOVxyNIgwv7LWLFRKLMqbji5jxWIwAaM1H
aOz2shmAHGZBep1ebN2pO0nu9MSzgpMXCyoLHCuZnqatU4nQ8PzOD48hxF9eTZ1j
2+EpF+uRVCmA/EuKEJcyjIYode5f/hcl592qiVIIZgjEbPudYJRRjDqHqmnd2Zox
dC7Ue+BewUkPWcGSmeRJUjr5Uu3szXZkxWHBpFqCJxf9Bq2V8cxVFUEobAwCwtNa
YIkyTs69K9ltKfeCThIUwKG+4i/USs0k3v6fH1SmE2h+GlnzH7uQBuWTPXLwuMmS
j7BRCrZ60k1TmA1T842Degln5JmmjQSBQHfI1R1En/9kmXISkD7BwSseZOSz0fS5
y1GDJ5ND/2SwFsI7m6htlc1oDRDT3AQedjWZuXr7WOZ+9NcUpuTRIp3mOo0yp451
OR3LkpmoCINIUuZj6qbLtvIwl5siP57VGT9k/AOSh/EYoJljPdp+b9FumdjQmPHL
IOf6+Z8a8x5B28ZRnjqy3VbdrLAA4NKeXOyVZxWGF2mm53wOpQYtp+lnslrhgyzm
qd3Nsqecbuk55qjWKXHIDms1fE8DMqjtnL+QBX4zTaN41PzKOfSvaNesWc7VhNAR
YNJgvjwYQeldTBYxypH5HOKPjRhGPH2HrOfpXfflrwO5MyBgmQXxd154k9hFD0+A
Xf7CBycNwMW/n3KBnfL6xcQ2x4AIRUdn5+sB0BLS1L4hlnH2w0poSujYIq2paYiK
zuSmMf17jigaZjc9bmLWEe1DrbGSW91lOeKrdrkz18dDxPCSxqE5Bd7DiM1TNyRX
Bz5+QIvZYM3ncTX8e/Uahy4bLFZdFD/ivOTYiPF/pZ3PzN0KaN67qdWowLldT1iK
AekJgaismPpAAPZn4qIRh2jce1DZuYDaE3XhWbd6M2X2Cdd6ZbDl46kAhdQWX8uX
U9cC2UJyRp4e58PA5XSzqWZsoag9mRbc98l4XvUuE9b1LZmSENQ0wm4+cvca2DD4
NLKZ1V3bpZl8EkdBAInzHgswqspBDwEbXSawrpVdTlMQ7FlpAk2FaFpxq11257rG
WXHDLI+RyKNe2PijktL8YWPOv5/eg2oS2UOAyXV6wAslASISu12gMgFgSbPMlsVz
KNaDkwdTJJDlTihEjCCWA2oNJl525I3+GNSexSRDEHaUpBJPO6iqyHcX93/2tfhb
JRN3aOGM8smUWZz/Zj/dhWa1ZNGXJNdaqTWo2ChUgawQHFPMQzZ3n2D+6wegjOKN
oWuuB2NJz+/TW47w4K8wkw4FmmTdB+HvwVu151/vt7fgSVltI0GUt2CKyExXypws
1/OArogd+0UlbJLeBLPk5iYSSbja+Je6plB4qEcg0FSWSH+oga/VVj7hxF4oNH4X
BS2hxqadaVOPtRbSdTeDjU+/fmrib0A4CUuWt3EPyudadzDWG5SJAk+6X3L1fNnD
j5TDdiM0oKrHRNVVGNWvLKLFo+pbK9sdZSqWxrf/A5bfcjVXfHiTatOUNqYI6Mdr
zgemmIp7rmM/I2l+N9mIQsUU05QLviRGxfZVHSeaQSmNR8JszRTsjX+wCLQIlCki
djkcFSUnN0D0MPADCvk4T/NHmviZ7EmYF9M+1Hw8mrGGXvNvaXXn/p5ZquNuCwnG
5JNPFwY8ob738Oz2/pfmztflLmUwCf7OvWjrk3p3xFt9f+HDLlztq35fnHLhHBXm
ZoYE8VWAZHhP0k7Z7vDI/KRYYG2GBQ0bzsssbUyx0RIVJtwKH+AxKpHNab5mHHiw
EA8DECKle6ZowP1ecFgKd4b/sdnrJAkJBSOIvcDi+PotWL2SMTFOIpZ7pvfJXA6b
DgTIW8X/RNM0AwZold7SL/o4I1sjaasgsrL7yIC+0WiNob9z/OnHBBJH5U4zK6ZT
ZjYtNRWImFG8E7Wjevrw1roNSCd5cHLyargwsLbadrPKPgwYzY4u+jSjFjLjZ9ip
RgejgX0otWkn2yN1nUtzXURT6ISuGk+RHSK8q7tx7wifJv0ZjEoD+KR2GBCDeLwY
xhumE/+ZTyiTDbe97EVrBqm8wveRbYHV1QXGp++zp0YpiClSQoWOjhXyyieyo4oS
wmzW25GzxEqM00p5jhwQSY94jKtZqMqUjO8VX3uPkUXHvvFbHRRIgi5ybjDFCuM8
mf6S1ttt/h+X23coEhwo8tbe1FIQQB4ccUqgcjv2PYLx6rl0ChRVBpM2lSGC0UnW
XaaasjqFIF+bLqKwGI0Nq4g6P6miyYYGlB/Dlh/TyeA1wZL1oDGdn+L9YgDF72/L
M+nfJ6JVqWINxO5YIUilyTccvN88Q7Rfu3mLfkB6quL7Uiih27uBj89Rl0w4q7Cv
YmmQ2gGF3W7UnzNQQJqPZhXrR+2b59jm0f5glGNnL58Xh4pnZUjLmwg5MftyXlzQ
HLWAoc6cx369e74ckoTeupG450OMZ5K9GmIhIHDY+wgqw0lLrt0rO++WXWW8i/u7
LbPVUUo80DTBaGZ8nC+hWwIrNQE4OrvCaM7ImU+nxj32CB7RU+JyUHw4tQBTH5F9
7sff38xUnR7KypANbmBV8MlzsoAfamefwWSKDhbeiXJ8huqg9RlV3YX1SUWQUxcL
DjEso7Tur6B00Pypd/iNjwZhx1FpSpCPWQsFEl8Hv2Bnn3ENo/ojDYC/WZ/QoH6g
0LMDSF5ZQrj01xFGsLDfqt4eAkuoS575ajQue+bVaRXmDyiNBtoBA3MomOdP5nUa
xSejqE6g6PWcQiT3R/v05lrbGkjoGMhK7ODGH8VsMHHf0VAZILsBiyCF9ONA/xm2
IkA5v6phQn0+3Hi9RUEk/QQjPl+42dipBZNyiZjliqw7IWx9TkNSmuWTHeOnUEIc
5wfpv0VjiloemTKAfoYVi4+gqmdu9ChHuleHIYIp7qn16V9EG2Lagt0VZUSJ8diW
AihRZc6GZJ7fTLOirjodB4PM93dZ5LV8XvS2WmyTQtI+QpxXnr6DhrXIUyp3klN6
A9T/ERJL7f6BpF/xTbEW0yeYhe0hbnSnyy54Zvc4t8o2h/h2DRAykBEp25UhUeAv
l0LXYurGxmTSbwKm9MjM/uMVAfyE68xG24ULZt0cu5R+zEYZ72jRNqmGi+dRaQiH
DKvs2gVAqd3bO5wPRt+AvPINsM5SeD5OHcJRbVb028XWkk/7YF4Ihaw3gbhif9wZ
9QHLMspCAXVjlWTNAYg7JnVDLEZvQI8wbcqj5C1lyYJHyOqPnrKNdldTIqwh86Se
s0NNkfEoBbgwt2mSzghcAYCs8knCynZtcQaRUJzUmG7k19haa6hBdBxD9F8TrSGR
utUAFFKCvGqUB6p7S59FwCvzPZwgXvpj011NDYXSovzhHa54MexEV73lkIK55RXT
QloK0sjCStWDV9wY42+822Z8psv4r4bELd9uzhN4bXPL77QIuRG7uEfWdTUnhMFm
NOaZq7ukf3W+ucXpbXtFe9BoLsVUMNwWvj/KOTsyYGS4K+JpUuq7OepvNlgwXPxc
eumaQiFU8cayT1fHsuthPzZK158hXT2ePYrWDHZJrSqhqMg6+CgWw+jW/kB9OEhd
6dC742RcM3yxmbZlQq4IKkJGPma2BtrchXopdqWMn6Czr9lmoFmzN+KAjUl+2JR4
MYjvFyTCvTVqE0IVA25cLunP427RZNe35ePL2d8igI43pn7nlIr56yd+Fk4dhWBL
8rfoYeOCMwL7ePyTOuvRA3/zmGnRq6dneA59ErHcP+vZOPzdVg2nVCBYsgeSQZgc
zxzA8UdvCM87KHeZ66jE0w3XmRAhoRxfESiHoJeNX8Cq7T1PTdyJwtA1o0TKwJXa
ZjevKIH0TAAffqWE9CQINKpPaY5/Y1QrKq3zUeXFO+JzYRTZObeHcE4+ZEvr5rbJ
1zzBKsA+qt3iLrEXccT8lV3FEXm0nqcJ9niBff6ZDGo2l8ZKvmtzaT7xJNS6JIfY
m26L2BhF6+yfBgUmOx3BvNvT+3btAO7Q893ABiuwcQUffdTUblrSKI1Z0gdyc9jw
L7CNf4UyV2WeR0EC8Hbcgn4QUjiI7RaeY98JsoKWWcOw9y3qt6Cwwnqvjy62kd+s
YRD5g4Wgwas1H2FLcX6tKahfH7DsV5PQV4yzj7bZdYk9tQnrLkGDd5MPVymQC2se
gv+NZIZbEf9dQtHEcVIYJj3ZHi412kcFEV3cZYR4cxMYoSdyUIyTM6Yx5NVwz+ef
pBnxdJhGw03iBpjHAt2DVeF1/3MEVACqJulQ/qeRDTgYubihPIkGSga9hxLxy3Il
7ij5TWnzOThr979TRHzT/+YKIvpuODHCn5zE30QqjzIkhC9m824j+ZcPwnvtP3RK
paHau0FgUJLEzplD59qoRufuSYNyyQWIPKFuBSInxEHC/NEYgEzwU9Cf2kVnf2cz
T53/8jCPF6pxVcKsncWTONg3Cpdt2pjkW1mD4nHbu9Jq7fWGn87BnFwz6QOkMtXH
qRJqcvJCfIw03qLGTjGEn5ITGFxI/qHdSPQHY8UvnlDQW66IAwmtGT7iDD90dSwB
mwIW/+4qkbg8yehSrZjEPp/xeLGfonrjT0pLBZnZQRbzKuhr3omovZtGFxO/PaTp
oxgL0RLzIggCkLZC1DXZKFbA8rTxq3JXv2DghlF87xAdHGBWPRRWZE8U6fUxJtqZ
PWxpEBWGiwpsHVUKTWV6Wdp5DHVXAYQCopQbUddTcqnBWdqDvplBBDdziU/XtVDK
mMgLehe1nkXt5m0rjecHWMnfNbYDbqXgM/o27LUTtqXLJyqYjdZY0LkUt5vJSt+o
RMOFaIGgCIRFthoNx8xjVLN6RZMjmnSG9PRgwsshSKNc6SbsycApFL+gL7EpqSU+
dqv39Y5XbsLbKM3EVZjfmzLbsd6biG3KRCZs6tii6eAqg1nIutm4CNpEwpDcmQUq
n97rRYrH5F/wvxLJgv+MHpP85VF5GsKrWEKjEZjJjDSk+I/xMZ4Ypg0wbtvazOrv
IbuJmq9PBbFe+0aFTL1bg9dv+ty2iPPV2Hxd0g83MV5JrOOlqdCLpXNv1Clqo2cK
6ipgMCuLnKM3pHTwqGTnvYkvmbByjuK8/zyvouAS0nPI8hfPvbkEHDeqjV6QNOVt
NK10/o7+X6tBJYDMd0JDJrQjSevd4M3PnWm1mGDW4pD0EdQAxUFOdJpeghsu/E6f
tpzyDmREfvlYwrwYRqwWk+2HiH7s2byB6839wUkbgiRFPJuqi1SEhXeBRnsoJafs
COoY2BHyINLLZVK9Wsr5hSY72uOKzeruRG3H77l2E3OxjBKUqYUKuSnwsHcgiMnh
V4pjp7u5K5NOkK2BRV34ErYYnHZ/YBnl5MUAzgkXpVwspnbHXR7zWiC1n2cTISXm
r3EjJ1aJ6zjf/PXgg50A0WQZbQARF3QNfHtZTWAQ4KbZKJyFxEhRVOLorPW9woIo
pNcyaZVoLcCGe62P9+5Hyq/litIlA8XRtG7DqbWqT4PUaunub1HGEqE8bfvjrxOs
aCu1PZLz+GqNikPgY33mefzlJha8uVzPJHaeqcbjHPUnHylpObkVBqSAWQ1CLhpx
9gHpDwAsKsxaXR3cjXOp+G5uHv1ELRhoyz5jW1qosfEnN50CedtX3Dm77LPCvrJs
VJY1nIRF6bH4iQ5MoHE282x9tHVg22saeqPxgA66s5iHDHR4EEpCkofvBX4k6Izy
S5SipdaDPIuaRKDoiQU6L9x8D2PsX9tidmHfHiQ7ssrEcwFOKFrw9y7mpQOMb3R+
V7YFrKrNXgMaMCiejeX3Uts0cnmnG1DR+vbvSa9cOWXKuujManxO3N63nGeQlsbx
vJ6akFQY6rCRywPnEBw/8Hdg8PB5IPmAckPu8adJPD/vwTMXfpZsxzbCynL2MdPn
1A8y07s/zLePCF3pmBURfXZ0mAX+eFJmbLqfqCB3Xo4gRoFaEdz7Ej423df50S9S
yH2XRk4IWDkAPrLt+eXmzB7eNridPwbKJBebKRA0ILXGQvkRhSPAbHSZTnnKSqJi
MPUPrwDGfyld48CaL+xFGxI30h+ev29BO8j+CWqBCR5M5nkevrCpwIOfj4nidv4Y
jYZcnwcw8pgrzlQQ2QExRCx1LWuwbUudZQS181s1vFX0xkHW6vFms1Vmhvo7h1CD
amadWQ01Q/dhUsUN93mR73atHBzbsqWR4F7bs1ITNe7qtivGw+ZS1l0qp4lKihHw
8YOf8RU1ND3bQzEFOVgczS9TfXcwbBjVpQJsruZW3MXJBvpcHwblxGsPKF4UN7e3
AnxNft0LqVeLfUutX3aq3T4Xj4tz/ZEV4rpXSMV2wIFRTLGQ+DiHFiIYDGnePaqm
F7YDSk5awbyK1og4U9Pa+AmwRhAcA5bxczvzICEOFbdf30IaeceC+FHxJcuMYWOK
r8bjTKY7QFGNsqoSfZHvfzu8k/7lsqq9vNV3vCbyh8rZc+XQAbE62F9fwlpKDaic
DhFplPNbFfPi/9CrCt9m9NgpIyUcEBuvxsdtd9/s5LwONYGuzMjVI43hm1gBC+k9
ANVJ0B/rx+AE+jApg6WVQuZ5uXEqV/x7a2FnQpIdA0wXEnhFk3tIiChit3+m7ovn
//SCkx2eMDImCiyzWvd898SDdUW0/EDwmCBdTz/LGXO869CBfvzFS+z548jnyzey
xrfO5QWqE7PofthCKC3Kxhxu2DgstB6AMSCjnDocNzmNA5na615IyHpTmDD1aN/M
58x81b8bCELk4/879w7y4flQMgyuhvVQmM1fM63JWHpGe73HGAfAPy6wpTsJJSUC
yVyqjHNdy6UX/b6zqFLUWl72tw5Z0HgIbkLrDqe+0HYa9+Wd+AmksZNCJ9+wkMeu
549MOlDjjzVok2nzWrDrrR9MciTLwTMW9+M3da4xs/UrouKzEyZrAXwb5m/5SX/n
Zm6cvBZKrKKxz9nj3S3hQO5PSJyHYyoFCzSFZyrgmG8uNUA/8f/1AVxNJLzKT74T
uaKdRSyznzQGYN7Nk7oUHog2G8meIyUZNyHRZo/tSUaU9nyqOthgqPl/GNNDatUq
8CTQiX4N6tKGluMQCLDkF45TO4IfN5SCvCCchcnoto2Y22ERMskZcwkqKWm2pEMd
ryeFd0k8n6Z6brb4WGjT956PZqsyCy3F6dKFkU54YHb8IY50eG+FvZfVfHKTzqLN
gDJ3xW+CWhcJQUu7X4huN63go3MzqUggTShM9PJuPGWByNxURkPNhO0DAm1QW/UL
O+xgiHK4tAkxN71pR1zmzSpVdF0C95xY3lp576jXJz1JdG0YwzkR1dlFtfYy68GF
zKQsYyQpNxNZy4MOtl9ZBXmdOGub1/dUqP/LXOpmNMO0eyNww7tsvSJJZ42QIOHh
ZrM4vwuBHGIRO4I3M9BnIzIZYWFAWUzOC4IQmU9DMwDuF9l4ygLY6XHIKI10HhMZ
3h7TKlLwMknJmPkUj/D+FuNkDBQcRfYdtg2YPxavlFx9YGlKuQwyw6ppIWO1mEVV
o/fBTkk6/9ndd9E+DyppCmBsYG+BNBSAlLdoMEzEb+eXast+wSIqQ+0WzDdC9FJR
1xpk8voph87m4X6uIZhRyU0a01YIc5RZN9j3AtINDg7JxwXywPgGzyx+0hyyluYJ
YIQnfVnwm6FDd+VKdihD2sjld0t1TF9vmjjdIqjss7hgi6S442rx+jF+OBbvXyad
CVtwDuv4ZILFA4bUbbeMCH1fnIEKoqYwTEYSrefotoqPuTda3Ftb/V4jUMUG0EY9
xCCtLpjdnZRW5WHAhB0hu8vn2IBmKonuRXj15ZM6jTvQFjXkQVWwt5p1ldUzr5N7
EmZiDk0trqKlvxvhUGp/CY8g9vGv+4apP0zHkY8+tsQjeCQJ4lDdlTt6xE3yxn3G
BztqMQ4TN0FCRRkNeanWLRJmHOBAjxn+SNMheE8AGhimi42hLtmT+a2vKFoRXvKp
9vR+J6VGm8CFzeOe4qnSFU/Y+GpAV/46dfOsy0qzFt9YuSA6WgzP6lE8c9HH+6b8
9g40suOTK0sFM0I5qBMV7eH/iyNAiGXBcYfnd//kLzFD+01c38ZlZ8nUaTCGE6xO
DQXK0gBMJ4uEw7+ev0nDkD9WkOEUfms7P13T3lfiInoF3ZPewGKXrQnm/ZTxO8eA
UhlPymaOVzgfuo6hFBnM6WE3BUrl92kOJkdOIrKLakAa5gLHouQ4qNFfwZCzBlNt
e9Aj0oyzmPdBFhrccSV2p6P34O6qYpKxQZ9yHMOjsefUIjqzQoZDlnz77MS0yvZr
RALUayu1E6+mTJOhb9OuXxlurf5e/D9dq4ONhgyCM5JQYge9nDZzRxLR5zEt4mRE
t/7ln3jW3M7v3EmIXzEEwiIgqCCf7yxtNTr7324d9BaiCDMrLYUrRzrwjhuZ8cdo
5o9Gobge2chaRqlXZjSlF1sfTZ2QuJLZEAsSG/lrWcGRpBGQLLoSNCojNda75gmm
vyBRsJjeA5e8DO84aS50/wOIpe/WhivlAOJ1goasJQxRUtTvs8vRtwnOfMVSha+q
tdYxPNyaohWQmadxlwYY7lMB2mxWcs6A/WS8seqzJya00l4PNO78U73Cs0MFiBt/
nHnhb6EnnBPjoqZHM+EksA6t0tD04YgY1tVLRZCtLNh4UMB+iZ0zT5O545A7upxy
0eeUB0N7G1kohhfvWNHzqP71HPtWrHYezsTXrCCQ6RqDycaV8v8bLOV2xaa9AyKv
oErvYYlq7aH3KBZSZ6IMcMa1kl+nw07rkvHFPSU0fVWwVNL/7+2VLieByC+4+SHE
rXJwMI1TuRW0zVBJ9c/Us+cVmi5kxHnHcEH8mxx1NmWcOzps6LY2K2XMH08/w9Pe
qkQ4MnfVdxGuGjXOxhmF+gv3odObA0CM3ij39T0hgQMNlqL7dDV9XbafEQEm3mCk
iChl3VOv6qVbutLRNb2OL1XzFVXcBjK17c86pT8To6KXBSJ12rcZ1oV3Ge7KKVZN
QMipFSOUlq/PZ9+6wxy7WdngS/nN2A9mkS6/WIIprco2REONYM5Se31Tdpt9xG/a
dqlT4lH1TWRcYVFIq0w+MbqnRldCz4UFC0PIh7EpgPEEEACOYcC63hMQ+HTOfAjn
miewj+D2APpJQKlse6V+CzjksAsukSlGDplme4+6jZlKg1F1nnAZfY+ojdxS8ZtT
SmcFpA9ELG680nx1yWPtaA3G8Un73nzqLvdvvIe43Rw/JWmQFMM9FBBqB2VtO6Te
TzQPII+QeHbkcVigtiDFpRtXWgrADQ6qC8yg9Jef6i2H6R9LG0eEN8sZf9eWtSD+
S0Woj7kdIcUqFMEUvy394bijkSs4/flBLbJvOBF+5CcLbUfAu0cVnkszIEDQAOSZ
sq9XGBymoRAPaFl95COBQa5vFwxKaK9+oikdBmycMlxkJhh1uBQVzbHnlJ9nubLJ
eHZZB9WLnwBB7Leg/q/RXcVA4KfUKaBEj69Vs8YoKCmvQwDHe8CXchfzuQx2N462
O9W+bt9bZcdyk17uRmtCgUr5h+rkbUrBINkoHOpq0NxufUqXyJXfQO4W8aBzdrU5
+rkwlFufC7b1Jk/do0iTmaeHN/b6XUsKwZO5+DP4I4xIKU0mLiTU6ng936+nG8tu
mvr9yDOOF8rdHh1j9Jk+5cdskP9kuy5ne2CZjrhi5TbbAWPOTlmWKDpZ2wEMSQoB
n/v4183B/awD+k7fYZtXIr4ThaF9mLdnvOcEle7jRrlT1w43/cbotZeF1OCQr0Ix
Fvb9dWW/l39HdX9eXC5cD7swXehmridATd3RC3ucCNxijWzKgJQgQGbWrG55rWXz
hShQb3Ujhe0JpoQb63R93CyxmJoeJKNemg8C/wjoiyUR7WEWap8chIwoxixQDPAK
NB6HdQ4lK2HEtxFU2QaUn/PqOdf69ICnNSzs5Gi/vdoSo7PDJoBZpe2iQa29owfA
A/xWsYg7liYLFlURPs4gTBidYjT4Wcrz4ulANkSkVIjhNsZTi9bYiSh09m3Zcp90
FHBPdGwBkD8moUMylaw6GUWXVzC39TgGCjSjF+AD9easZM0Q7BS9WfgjTjjsMqng
VnXrb0h2qU3yLVwjXiPdG9DseF25Ad8Eh5hZCA49ZwcCNFD+pGcyrf2yogoGz78P
wsR1F+SLXHnvfo5vpmaToYYF5K/f2kSSHHYnlJdBLCwUi7qbQtol53I9uaNSZQQk
g1jVYHpaEHfSOvvuz6p46c7PNy+U0csU7L1X4wsWlPsrmzhpKLMczfSoH7QRCGgI
e7KNj6Jh4lXjB+/TShjlG0c8prmIpNX8Enf08SbG6nQKQEWPSNYNwzNfNf/6w4eb
VusuGIur6h9gpocfBNIW2IAxQ95R0Ot1VYmDfcXmXEYT+XvvIXEIT6MFHiuoGHOc
hlcnJokvMAZrjHqhticjcsCUkqYZ6yB3qrbdyPOaW41C+InOLKz6OdveQ6BSPgjM
rFBqEuxFO5rtHchCi490vapruRy7tW4vnkj0v4uhAGaEk4xGMhCF9Gm6Tl8qFP2O
+2R6f5MqEoD5ef0Ki5ag6t6H0i9AziY1w4uqu3XozhN97QyocFeVG+yjR86dgvF6
b3Z+Pnu1e/YU5KIKJWdTW72T0d1cRUZ0svvZJxq/H4bN8KCUr3HpOKSQwGsl/I0E
XEcF/L/0PvuvQdl4pBaV81KlgQaisGSFrzVn/9Lxgiz5V1jrE4IhdVcoRU8o3sL5
/6ls9ZdpQv69L9GJoT1mQkoOr2VfMHAUhYGudLAJGTApi/shk1OVAF94fAGXEa0m
rVbOPAT4clAIt7I8/qrD87sdoZgVlclhgbQMAyBnk8SZZchoobzfKNg9KscX5Kw+
rfaTsRaxqMNbXT/Dl2gPwFQva4MFH0tVCGbZMZL1UdCV/3q7UhY4Uc3kh0NOAJdG
jYgl5loIKqzk1k5cgRsY53wY321fVtAHd9WAE3cwpi1EA1DdBpZk+T0h/vtF59k7
zsl9YXrY7nr95mY3SAJgLKZcOtOK0CN/4XQqkgG9V5ylo3qhNs4spXCZ+foJTovc
Gch5HHWXBl4gRp5LDCVv4UhgiMRNRbUsBI9MOYzqLhPIilH5dEfMqQ1A536cffFS
4ut65mqsUIhI6lZo2TtlZ3NJnKEXiXjnMp97eMouy3RnBssb6f40mv8FOqszALX7
NU63Typ1/ABYOq9XHmpzioxMKrtj3kRgRnAMpowb2/SbKMCN9n3OK/kQbUzLijwR
85nz/cRGiLwwSy8BtQxZr/ztEGpsXtPf1gHax05Pu6aubtUNuL3b9QtVw9sdOKCf
3netlFXN7eABwQ33uOIzq9uc/DyAy1P17IHFKZ7WrSRnsKjn5VMRu1xsOO23hamE
mlT8/+BuDKGBW/NYDduV+VQmqa2A/vJbIopglif16AdadV5dWQeCPX/Id8k2Kbjs
0XsqgTdvQ7K9nSLPtOxIyO//Rj30YlM2tNaKSYO2PNWF+Tmt+flYB10nI9sKKvIA
jicgZrvSFZlMFdy9C80zCtJS9dZytwyacb+B8S5/QH3S+MKQbvijgf0LofgDKaVv
s+8OcEjg3bZbs06p4gN1oz4t9QthXaTvdEHV5SG/X7xsi4sxTb/84jOACae6tHGA
IKsj0+sv1brWPPIjTyhtT/X+brFjjCsgaF+CCud3H22PvHKlVzFneVzxqyIZZt9C
6U4CmxkHESSe9ek24ZNkdQoPAr56bKcy+/X/OLkvsVh8DGzTKW8NqvV6N7aj4QqK
tyDHlWvCOgbz7UTXz9Xs7acLWyStP3ncJmRsI91aPt/xkpBfJ62Kmr8AW95wF9ER
Ldy8A8LUYSxk82GIe6Tr0xxEbx/34L6SOinVTC/Eqz6uWIuCVAtMYGYREMTo3oK+
ECne0HP4H/b+z9NUA7sa/akcFhSSlYRV273dkf2aZTZnuQgE3JPl/TJt570Wojzj
UC1+V0NYu7zXYhNi7SGAX/ME5YU6/MS/xWBNSSm1F3Cj+O5YfhXLLuh6suDvLYh9
ZpRb91wkjqXv6CGsM33UVQMv4/T1Nj5hGDOWqZeqlrWkS6oheNpFXcT/LxJ/QirX
aXSNUsndb8S1kvWJVj0EWB+VBIuMa7d5oFsftKXLv/vmAd/DG5jvW81b7+KfZNRw
mYoTvCNr5aSHy7jmh6sJ6wJSO0OGR7wUaoPuvQ09ZRBhsX4DOe1m5NBRqgf0xSlV
iMVR8Z9pgts/ftOxjfW1RPE/5sCPWp5pue9cMRsQMmcmoz2hA4zZybcEj0B0ZPAf
38L0pYswAXJ1oqANuoJzHPhBdVr77rliYmsldyuZp+X6ed2fvjBfiyZ6xeecBY4w
rWJ1hG3wrjycW/9su288TQ1te3qAi45gXySVnf58FyKDz7GJ9zybjlmhE1W5x3hQ
6AnpuMBuz2jX5k4jcc2yUSW0sV+k/JMwoUtmrfXd3Jmaw6EPj4fOA7ZWX2KyVDQq
cnIvSw9HCg+21aYCQ4qO6gVFA2QzA359wZ5V7c/lBK198BZODpdLbDsdvsfaeRG/
uK7eX6zYtyw6JjEn/NtUt3EuwA6sfLOonQm0CvQ/ZbSNlx51hQsRdFU1G8YrEhbV
QZcto081+6Zafgh8tvBKV6d67NejjUCqhgHWEQ2g5kToB7wPrS9tF/WCaf2lNCJ/
w+Y3qlQl2a+EOq/EpYGKsWctVLJYYZ7nX2wTqm+U4mmKyCr3/OeS7DNCll8lqHCJ
Z2sQtpP3ImcYvpq13emp6+r36TRByURyFhx2HgO/qaKTWm1nPVvRs9FGn/5G0ump
5HA+UchFSBMEyNFBnFmTHphqZY1IFk33tahu0wxKvt5BFtGMuxidYhhw4pRgufFZ
BR/7gKD527fx6MzWbp7PXXUMnN88f2jeZcQv9orqBAl8lqpxCzwrvZg3EO4C5rKY
4DCtq5ax3ocZAMukdc2/O3FhOv57gdTfTuntJy2iVOI9Mm1lzgrT7Rk19oQG12x2
xY5NxnluFDDcPexNbTEfgL8Sres7gRppRACrtdcou+k4SaKB9VtvERbVefupUPSj
JONPpGb9UZcerYsYuvC2CdkwSVh6WXtXX4sHFDiEl+iul4LAA16Iu/ZVnWV4iFiU
vcZpCXld7S/JD0i91fCxBWFRX9y0J+dVIvPEklry/kPQt/R2fU/2PfEy3DLaYnm9
9IwDwSevIp2ULFs2IcZx9NJHKNdaVTd/LakjKg+IfBFW1CU0NiF9J54lXHHiSfJF
PLuS+rMXZ+pib2WucDRHyQHs+yJAvGBkNgSj6nlX34iLMzxWg0OZ3vZmVphT3PjQ
F5xazqTiekZBE4/48jAZ17VehpiuTMruVgz63L1jofqE8at6FJmLM6fsXJVGU0Iv
ZP/VGmUq9R2JZTCIl0ZQukDR5I07JEL2QzI/KzJuMKXnisJZMMAK3DUd1AHOce3m
IOMeYpzlDMBixrg+JCVrQck5rdae72iE+gZ945Y8u8m6y/KWBteHNBEQxgFk5eJO
aKuY2Yixw4zWhBMjeMGsFNblho356+wjO8HKJbvQX9QrSArA2x/iHqR3RW2NvYPi
lKzhhLBfPq+ZZF1Zht1oDCYiyfTOwHBqVeJwnK4fkIUBUdAV334MkBSlmV55nEx+
9jUjHAvpMwm8gb9doRUz1+ajMCK9TsKuVQ/iuFTqmAw0NHehT9wW9nGQozuubfX6
HXMt+6NUeuP4poIto7YFCDKem8R1mFB4WcvCXx8fjOn/Ce3msMqh+53u0JFNfnZC
LWn1TJfl6PdURBn3ZwiwtSxDs2Ijt0/Q+IoPLeOGSiSGAUdOaW3ZGvPzCvRMopKZ
CTPIdkQhBZgCoM9/15zkzSEBGtqZuExK+gqmPzrFoiMTwnUjWeFANHtArFoZ6v46
sCJLZx4SNGhPQ1SH4emdYGdtDIEwjw8zf7MgD3lR7oHrvbZr9hAz16FvlqIemxsp
0122eAhJ4nYKsDh/7G+rcGBJnAVSZ1q0nBcWOGdfuSVxGrhlvG3rmXPmO7EuZX2e
aTka/q3Pot0RnOylWbePESnDJc0yD641JDGiYHXjENP6fLeVbzBMH31hujLmR2xF
LUbI16fvC6xGk9tNynal2qNj7dBBYZkyxeh+tJrHQFnidn3fX3vwSISoG/tWHpUR
FjetZuOq3U6oJud0XQhtwFgxVktMJ2ifuBTg+WWMvvltXjJScJB4vDytwl35TYba
AR7DPV0iL75/flRnS/X30I0y/HV5nV+L2/DIMLBFSjo5MgHqghbYHbFUdgNYo7Hh
R8OXM1bs1T6PSZ75F4mvBQD52ShAEtJz7S8GldUHL9ef+NM8DljA5JksAQhNwZLz
OidqQmhdk0fAera4MdkUoZTiXQgCP4z9cNZHLm7q14246BntbgI4CUupw+InU0WT
TbOELijsZXHQNHrpE6xOc8gjvbhLD1D5rib5/7EdcfuaiWIfA7a2UBwG8VAetqUG
5PUJCViBjBB3aZ+f57yH5uxnsx+kX2fhhKmmK4vJcB4FwCCJYqmYuP95bNNUywN2
ezKKsMJDsQ3rH2XWSDMmqKXEjWOBgbh3G1mg3bB90tFWDI1aPBxILeHabJD+Km0A
MjwclDtrfTnIahnFt3DUaFGKgkaq1EfQt+tK7MIm+ypI7MSqeW6LyRreCx5fscsN
KQexFlBzdKm4LPVKYfN1OeJRf6R8v9EqeVoIe8TIiRRqsHXKTMOMWZU+rFlWMd1R
7fv98/fhRBHSN9iJ3XYPQnP9kDrQcJy1soWovyFacrltp0CV34BRwn+hnx8SuYt8
CFK/ay1iq8gdTmFaOx/jzT5lXhnON2xmFz/CFhrUtMheNv/3iHwB8JxfAac15daY
9Z/uSj8oxWDo5L/WyoAhYoy0H/bBdHzDF2hIZ3LLSYy+L9dxNTMQQSlDYyYaA61h
sBgRkOO2IHqhc+5enODBIltpdIOJhuXC/8G117tqomFTGta8v0++uf95r/yuGzAl
Z90yWIl3zxjcyncawvHIbGCGeyWVaLV6Z2JaF+YUl+NyL9600d/rrMaSVf2kl3Wt
Wr2/KAuW+8kIHikRINgx4sTHuwlwe/PZWAunVDl2+eUC7XmbduX7MbgPnsxEADbl
YlcaGxOmGgpIO0j2YhGtKMfo9o1PKGY3YDomhfGByau8Cvhrbyf3RM4lQIS7AyZU
QlXJ/1V+42KDopnXnsRTJyd7aW5+knrEiOEz48fVoRxFXg73+ShV1SF4oi0WUeat
+pSrvVRkQ4h35nJ+esGLtYOmNyt02GcDOnBUOXLS1Oqf/WMc9OC8RaS+TNW+Y2y8
uWL2vKSaI/ckdtEGniKRXs2N4HGYF44/NQYBaN5J9JoHxHqcRjtbnU+IlGpUYohG
dyHI6BmSbxxT4V/ug7HLKso/i4v202Bm0SeETvN/978ggiNCUYSt6OlX/ChMhcaN
lI+5+8PQArLbrqxfEm1+9c9L57a8/lk0anVezMRTy7u+1wQ3Jig0lq1kwElVzKkd
NYl6PFCfMgGPcXZ2rusRni4MQB6Eut6M7/Y7H1CLAtQ+qsURQLTZ3THu7bnB22zU
R2Ox+6TrRYTOTM9T/s/wv15pf+98/b51dubuB5erBpNh/RbkFFGA91MAvwefqhgK
GJHIVl9PMEU2jwHG7x3XmetUgRro6MU1zZRCWQaBG7MX6ziYy3WEb9hmxBKlCN7W
sxjKZI83L6dMyWQighkhYkGD4l06nK5O47I9AtiJRSuiIs+LDTD8tiaDr2w/Chig
byebcT1zRMo0Kn8a/9WwAixrdU5eruCBkjMAlNnEFX9VoBJLT37HNSBgve9LtJ+9
bjWsg2aPpzGV2HtmOqu9h+Bc4hpqJ6VjKtesYTx8u31/DKMjguiqfp8jwurI7kHb
VaSnpDM2A4+/Np/8Sh/zrDqm5LAXsiKBEApPnVFWAignTbmBLNAVSU0qEYv0NNad
bK82ttHySRg1S4js8AkmJMHpFKsBvURvSdU1eBDVAQ86ld72/0GEW4opYkd3QZz1
zcSmWTL3HwDCWBLudWzd/nDb+SKxdRIkhzrPw2zBkv07Q0ssg7Wivivko9C0oLju
NQWPS4a4saDbm9dL01tW4yf12HyV2RwLK6DvukLjg8R+GHCgDG3m4B/rl6n4H2Pl
jXVRdoGcuKAmcbefqYkIJm1tIQwbzjf+e4IdlVB7hKu5M2Pg+1Q/Bcn0kWYng1lr
q5SP9Ok52MFLp2rSDwT+07sXAg04FXZYPNz3cGIx1GlgnoYxGWrfLCUWnqjEKua4
ZNJl+cnUHOgnHMXjhRcS4BTej251LRdlWFP5zSdlHcFguQyKwND9MzG1lW3Ciy7o
tH3HEKu+2U/eApk2R+TorOybDJqcj30/l4b34ngERh2/yuKosvZGEB72NSC+ValD
4KPCgyDQm1Lkc+M+TnqIb8fn7LANlnPD1typsXTRaeT1hxGHGdGk67ubAZBTXEYE
H8ZVAGonWbTyom7l3fdxSolM9OWzkJNkvol9fSATupzdNY3o/Gf9zC6O/MSAfZSB
fx9kw1BtuWi9K36uWAvlny5lwiocFOdDWK9BqXqXwaSIY3uvToEuXbjpF4cYSWxk
fG98JVDL6BJLqLGrFWzduOIorZCjMsERoi4PrgKe1ePa63pvdUy+O+59zBXAE05o
rJ5VI0zOmuZUaV5XFZPBIlF0wNf5eznJ5xKbWbNNkqJanQGGh9kSCdVbVkr5wCqi
W6dNEVSBehb8OMsG4zOK22LPIee6Rg8Xq2ICEsxXPi/uH56sRLqtCuWNudkEANCB
WFCmee0BmrouNJKz7cULPbgSSrCbxMGrD/7Li7sLEITEG+E0b7vxBA4ORI8r67lx
hRD+zAonUxDOs9vYRkXIMKvWe/Nh99ZGT+SS2KWVgA3un3wc1vD+2fNodwk3R3yM
9RjHujnWjZSGyXZRn6vFHc0g3ynwIuRbzYISIjX/68mYx+BbjxhtPvOCtARKZtPM
b2QXtVQxNJoy5IoB7STFCVEucNLq1fsjuMENhawsMYvoZwUtQCgkq9qk+1DBBYA7
QRmzTdVrnSqr4Np0a3Yszma5bJBXpUIA68/I8eVak3MJdrmaNtiT1ZKPUGm+b/9W
r0IcCF5+Tw4OGmasTB8BlwqPknCOq1/afOy/fhonCDci09CqsqYDagd467J17LkD
Io2OqzlcpBBOZdQRIRYpVGsOjzqI/FghXVe5hqdL5IkmxHw7XAJtnbTC0c16mlKs
fLaCUt9Bj4dAOVWtMA01Eb1Nm8cHKhzkG8XeXGlnTm5n+YYYSV0HyTwYGbFh5Oti
yaQNoXNDVP9jP6CEFmO8+jNyjyEIOCbrGB1G1mN/5++8mN8D/fMluweh+uBuSjSL
oPb8WK6GObhTlpNmO06SX5LjhuNXzkKv2JTSLexGUxoBwbx4tob/nSrhDuUPLUR6
BzOpWRuQjcOcsK4HL4LC7tO8Ks0EFY1W10fmAH9pjwgHTX9Ti17l/JppIUx1NvBB
j1oOTJXK4LZyMxCtgsYxIvzpsqtCEZDdEOQcFY2GLSrVJ3WB2ou20fDpwiQ01sNc
2WHJv7+gbRm6F9H8UvgwXyMpj1CChD13nZWJ1bdXuABJOcyEGpyQ/3qiIPgxkNgY
FRtTJ8mALnZ6KmZIVoRK4CzJQ3nycXAEWYZzb228hzDXampYOVat3xlAOIXXIfvX
T47QtjKbIqmKUiNVX4pI2fjxUNNstngJcS6TfxcgK+4Le8vO+IyhIOHyuUTVzVeN
Ym1e5RpNlij1pDIvUGz/0985aVBev03tnurLA72XDg+MtPWY+OUcTuK+0C1HxAWx
nX5EFfRI98qFD7/mgs9hDfklPF3F8OevNZ6IMLnxDiia2QmPF9zpQhZuHyeoVnwf
3bHuO1FqnVL/9ro9XsSMFo9J6PZksjJOiw1F9Dy9s9dIdR9eiqogEkU5VkiEDvmC
2MsaNLGPm7QQLbiivXmYZTPCcLfzGreYEqHpBtzLzr6JqvrLFPirsKckE+fHwApZ
uN+So6K0FQsBrp2vWC3fXd1oCL+rPwwYA/SHbWjdFsCDMo7dBU2fh1tXphGGV/9X
Rh/8kA8JeROaoL9URZnW0s6vG0q4tjMPdwKbfBxxjF7woA8jT+b4ZlWovNz3EJSy
QuoFOZ6y69sRzdjZqptwV5V9rZTJC5XqEjwwAv5YMIw2+UjeiVHCdFlCr7sPVQTJ
8LnZeB15QO46bAWpA9rRvlYdgDq7XlTlbJ44Z+E3A/bJ5+PAt/Y6/BlWPBGRE+PC
97B/HxQGWfPdcfbpsJ77iACSs216NbKLVAWI41EPNzxabOpDDg5p/suwDtCaP4q8
wvPxcdH74Id6AVFHF1UbL0faWVl2dBsQAvMbVZA8Wx32IRFvQ1oQSfwmszP71nkc
fiB29wxQ36MgqtDMD1GjdqLiNKVsugq41jjXH1KG9SkTf/cuNw1c9CMXJTA0a/01
l3hoa0fU7CTpe5T+ELtuFKTQfzUrcBTwtGnpR8Dh75EvbkrCk9LO8h5yilgGTSSE
2qLcdq8jupOxgWwo9eUCIYXlHmt8N1mP150bIvsiwsgpBvbTrRiZ1GcfXUiLB4Hw
7PJ8ehp68CjMJX2KCAkpLuepvTGr8L2RkVUrTdUH5xWbeaxCVra2Qp0RBD0ROD9X
okqubrV02FX4Svfycl1h9qss2ExqJHj2t/IFHNTm9jiHqQK/w8w29cOzrqYjM/ID
wG7WQSvhcy7jIKpXqDazh5tiuPs5MqNGWNhSUAK8SH1wp5e+CJ157RSk0fzAonbp
ifu8l18z51rA8Q5f6swrkSxaHlkyo/USsDOYKvVQciqJaXMmc0LWjk4Ai5O0+zxp
+9KujCmVwoMAqRjws3LX2Kc7m5Ov6a3RPajGfUEjeKwiTrzsMjwucukh0L1JQCK9
49trUS4G2S0w3ON30+uEzC+V+1CKdvr/8p1AlW6SZgfEYNa9CBCp43R7PYjQMuCz
US1YCUGk4vN5nHkg2Xm3FW6x8inbqm1F7CNenN4Em/Ut/NCJ+RUGEzXsKeC+BP5k
4kB5r/ye5Sur65RxT0uQHIjolaDelJ2B4v4EHdZZMnC7jdA6zqqHGysrZ3RGtMu7
qOGc+i6Nm1veKLufEXeg4i83m7BACH/a3Fyryj4JnNTD4BnsrUrCQGzZ1qBP4zYQ
jumazs7xrAGehC7mfoqnQToIrlDQDpIXotUuO/OZHahvWUPohQr1lMTtozrXJdaG
9lfvGsqfHgsiEAkpz4JMejaQ45t3mHc+/tZ/9U9cMToZPcIt1JHMOAavpz/D0XUU
sAwtw6A73LBn/6ZeZQtWUk8W0Jrl2Q/r4w7ge/PX/SUr7h0tdWB5QXBtmx2FpyFo
FmmDJrumr3Nl2HRw7qnvnkvk7P0iHQFE9BfP4pA1wRe127zt7dH2sgQDFeLV947g
HrwqKowiwymX+bTa//Q05S33A4rufEyoqxqHjxUKXNBxZ4So2j7ogYlpsFGVRZYq
s8xhuiLg2PKwH+JcZU/modDCdDlz4SvO01BVlRsMw3WH4XY1sruJ0dICogU++ucd
cOyrKWNN4BfLI0HsoZPZA5I0sOhDRw7xVnbJD+7xakAB8WwaLnX6OmFzxbZJqPbR
4gTmUUvql7dAL1uTpqfKLe3F3qmJ3X6osCjBNM8qsXkG8WortD3UrQAXY79qjyO5
DHnB5DXhXnXQCJHkYmzESZBzLQ7JKI7zB1uM64sVE6rUVD3YRrf6bdHQfSRST4cC
UdZ3a8lCCbwfR1r7gVylf4PpVwz93px8U+lwO9Cqw1A8koWDky6V9j/FYfRyoUgP
zBN7Hbx1kPgL+V1jVbKhiYk08HdOHnOfhV8zsSnoNrr7AfAkCLSBVVHHRkazj/E+
N9eauwqB7u8aDgDHkrkbZx3HpaCfS60yzG8lktExiRCb/N0B/ACHBZ4mhQszLKxn
U+tsYA/VD80R/EK+jskWoichEvdVfydsfundJeq+sMPfJZ3lk7408sgI/31wu0DJ
2HkZ0QN1ykwk3uQoycyGGjC41XiuliciqrK2BIVOGpeuaX+JpLHTFFTqf757fPda
paD5WNYoO7upXTes8819auz8vV1ts/WsTMMM9tqPQ+aaNiA4bUOSj8mFWRSxG/Fu
MKled3eK3T2p+syRU+YCpzO57gZRPwHNvILzcqgD1PppifAegNY3HRkb9Cpnx4o7
9weEBjX8SEj6GxYw0i+GAm059Pm+LkDip7yM1ap4zhoudyfzOcZq3TnZgzmE/Dnv
+Q4BeesLaN7b7Cg4Rpl3oyymv2pT/+zRzFWpYz8pmdSXDrQNScKppF3Js9Sq6dsR
nclLLah4dHwbIAUS6GfVCxVM/k82vAlGUq3NrwgQspn60hBfXEyPEFhpWQ/2ahsa
OjQanZY6WeYNWhLXm+0lVeYVMK8b7CdJSrXFseu49gGC5tdt1ZC5hV0lThOtc8Fd
a+9WTR8yu2HDMU4fwzZ01629pZ5w9dTHWL/jvAkv70Jvs5XVgifLf/8e7/3a5kQ7
+C4bme6Ar6OejeuIlDUeZ59i1q4W42FCtx07QYlSXMB+GBVj/UVgK4KaLMmu6dE9
eUZcO1EX7/7sAw9ww/FU8eXo5q08bumh2LYM4zki1RL2n3Xkxv5aqEvap8X+vVOl
6d9lcCA/Y2lY8y2mdgQif0MZqCMNYoBx570WqNPhZGfOBhYlPc7jl3d7saIIGDGx
SbYyyHP/8Vktquq+dxMPp5idT2sS6hprhfNZRATSaPzOOB+8rodId5Bxl9LeQrre
J/fth6LZHS1LoHjSGiW5gTtl4LxY7HWQ1xHs+kUAdHA5e+yyI7j6/UJjjJMSJ/uR
s9UoqyxK/lxfgqFwA4q5DWHWXNV7N5cjvger1TVqSfDG5+h1T1B9mV75Lm8rU6wh
u0Ri6BMtyNEpeJvFG1SRNuek1SYkVE64wSGL6KKWp+ZoWZzWOEVFmvZHKiyT1aNN
oOlgOjkS7zwT3rH9+rUagCxAwrE8JsaLzj5wiSHYtMcECltclyqHVF9+v/LIlRP6
zvCa56o8UP5aZRm+cXeNeXUioWGtqJBhOzagjXsz/3waJWNd1JTuOXiOXr+uqhiR
BuKGaUOckO7/oXvazfadOUmS/i257mZiNLHKyEvCtctqT5imyUT/iJNU16MCmp0R
IVCj+sXjFlzIq4itfxtMmSZkWpsH/01UyhoMR0xK1leSFcyGKP1RhWpMZ3sz/ha7
uESd7xILlLv2Tn2+P4o18UQS9I2+W1zLxQENV9a4n1xfyuQhFBry0p6SFUdxKkHT
feKkws9IhgtBovUAx89w+M8pWErFRQtEM5zJRfq16inTIb+unQaUe3BHBRSH5yyc
5aVX0upuks6l1z2ioLyWjpbWugYGi520SEjti4KLOr8WiFeveXSMAMsqQRMUwaBX
P1C/R/Au0CabaTjeywjbqG2tERtKKEPwGJQEYb4Gxm5X2lHRk6S/LpUux6S/iS/Y
A4nvALI3hYE1EnmcrYwQwwav0hEkfvbbtj0keIJtqgfYp6Enh1ZbiEQMEhraWHXj
p/DYm0aOF6Gs+TEzf669fJt+itAnAMyFypokVw5YEoftQYYXLSnXCUbPhsgMKi9P
FcG/qVjS7LQLlurrPJe18EmqIsmoiEtS1cjIWk7RTc4wJ6Bejq3+Txe1m2YDM4Vr
o4GEg5ifk+BitMgd63+7Es5R5UfVRj6vhdc3P5s8rUEbzO5EzeBKTsUJuBM6MgXh
iZUVOIT4+Xok1LvNmAtHPW295yo41S8CjHJAOh68IvKqK3wfi4y3ABW3UTP0G5RJ
wA7LMbLm79GAdh5/V1wIfFAhS4W7LJdnzFP1s11o2OXFNYXBQf4W5jPvFaYwUQv/
G6oBkkLWhK4V3Wv/OMwiKSMRM3Nr1EdTeboFlvbzJil5O3c0bd7+QixGY31A3Jhu
0+ZY+sng/8n3yV8o4Ix1rpCyNaJ1ahSWBuagIWCMkSEFGbqdqCSV+Ugm2LHQ9gah
ONDvTuvqCte+UyR6Qla08yYo5/lIpbfeOt0XOhtw2WLvkgtgrGU21GIRm6BElZRk
MIZYc4/zdksM8RAyqs6ZFniAiLi94VW5wj0KxVHW2DfBJKkAwj6yfHtII/s9tasx
THtvfKGzyx0UCMdkBpw46ZNkUSha0IJfRZfkxfk0chCGTQeqBvDnk6x5I9y3zKyO
jhF+nW1ux46bBoxvCIjsG+yj9LF6AKtDKQI15HbPbyECxOFSAsOTYmDDM/kxNei+
EORHH52Rok3noqtFUshYnhnsHGeEbH7OP4qsoVDYGNx/13EJcsIFAiwM8V1Svdk2
fas4RywSG6c5o5/zJqNz2pXPfDS1RO43Vw0M1ZbwOCOktCHtuHnWcT41Xsu6djwB
DDX5XjCJgjjxXC24NHz7VlUtAOlwulH7ydg1wZtnZMWDb4d+n0NSMsLzNRm6EozI
xqEgFGc6p2T3rxZ0uNJ0tu7XlknehcZ9Z5dhSe2eqzbB+QiCdP7EXlh87oNJM3nQ
8SFac8xl0HcgSsoBAcdwmcFv1jwUqlj3pi8ZmhDcfzhsUUzEy6gRpHL7Xg9dtFhB
IW+hxKE7dypqTz/gs0ma+BdoPnITto+NxisxA6lMLIGJQGOTtazpq0pQClPG7Fgj
bsCg9FLGlXHGDaTjp60cnJnMuKGxaxmVxgdorzHNl7RJFKUCY2f6uKqLCHEIwKho
4DZ7P8BdOss1t002kMFvXkd7wlvF57HBM5bO7kaSowgXYM7d7auyCbH3EDXPxu1D
Slp8gI/OLpLJIq68AFBjKJeJ5JTYyUxn1HYfbtjnf0rBkSG9BOS92QM+dlMnJWpa
7IYEytGXHrMhK+Veus3/ZAWYYmjygUkkMjpTnedpRSg0mhOuH26lfE6M7pAxVJH3
piamq/359x5rTKbmgXvH7ajgCR3YvhaLzMw5KwnDkB3aWx37IhDoPaNo0/utHSCJ
00AcPhu8iJlETsWdJR56HNyntSSqaILc/CSIbPuEFtShRSRpRtgdIB1cr+dW7pzn
+WSOVy1WvBr1p7pcmpqRmr+wHBDrI2tzY1YVFe6D5mUlNSD4QgM1bNIQuCkaVgXR
T17Aj9kj8sPAOcVam7Wy9MijpwIU7Z3fWv3ZRx1nhAo2Qn3RRYHtrKOhFcTGIJdi
hPpRnufczTTOgp/fiEPiafGkXRr96EXDjgan0C5Dy56tW82n38TT7/xIxiqxuhN3
nD4nA9pm7J4GFj3+EktYP3SFBlwaVrCAzg1pc7aydtSR6cgC5hvQjOU+ifAUfIBt
GlPGl9NVP4UThq9RGMuo09zRn+8lIcNZTrHIc8DQqYuIs8HJlVLdoXC+MDgnH9zr
32ilRuHibNOuDUT1+CU/3ZWknl6dUGd2dL4k0zLkNCHtEN+r7zeXa6AEIxwBWg/7
wMsvPBY5OA6BgyQh4UrF1ANKbld+ywSaCA1QVLVpt+ery0ZkaLcMNyCdbcsgjltF
Vw2r04ICGLwqlay2wcQb9/o213ERHQeieHkuzynYmMXQ82RrZEY8ko2lI60zZU+4
BNx2Fe2P9LGoI1vsJTj0G+Bb1XhLWozz/8MMWDExWrwNRqesJjBqZa/T4TpX2Wxc
XTtWUKOcxugj5iZU91uCFD+I7upFXj6SrrWrJMLifSSL0AMKVErebiRl6ZuFOLUa
k+LYFfw1IJhFXqKYOL9zo6E80W7EcD4/ATIgyW+S5eD+uy87iaPzyM5Pi5X3dOkH
dknSLjRKYbKgsEB6moOFuEXgJ/WELy/ylaSeTXVXfWcvzsaU9KeJet2SNRXEDexX
BIOrHrtd+6bPuEU3PaYTyBJGNWRATPGr6kDkiVvS5R1szzHJtTxnj7AAzlSQeAry
2f+S7Z6dkTnKB3JkJ10BZGo6eAMDpvj16PJw/Ar1fMJdh9EeR+4SlKY65qN8VgdR
34iSTQB2mcE14Rx5vaDH2nR+lPsMHlmsC5qgWgwXuT6wlMGQi6ukq0BO6fdHIX1o
7+CsduYKqLRuu6b1eFaFzma3nEMm7SypweVcfVYhHe8xA8I28RwRmbojahxPP/Rs
FCtSmiZlZ8CxI0H8bn+aaw2OcfTmkb0GNX3Ywoizg1PTzGuz6V3oMIqM69RmGMfD
tvhMzsSYo4XBXVJPrUVp8ADt9iNen0d1KnW2Ydrb/0tYSPZ2oDD4ws0a3+nknT84
Qsi5dG4pQ1yyBKjzaeBDtHvtnzFRlRtoCS7pTU6APOPfi4Ju5N5oKHjbMj8nFOuf
cwVjt71YdOw6cteL1gNJckOFmZcH2EofgnSCoTDGsGIVOLMepYT7b+UMaBeYivrB
HKxekeexJ0ff01sBPzpGBqqtQe9GZk6ovcUvJ9TQInTOZXumIBmogU4r8aJvSJLz
PoAyeVIFTZpWc0YEabjjPpps/GJimB3YErlqPryMrs0MMAOqhooH5ew9SkUUOjZ1
LnG4Zl4PyvcN6T2I/t8pNjgyGUO1AQsegdWCrb6JzFqzy8rhsUI82bBZXG0qbMWG
C8Qyzw6ALMepKrAQr5VmXvCRA/jTMQugM6hdK05e21gORZ1H6u5UghNdwcOuZ5Lp
cKrOiTjAl4hNoitmSJx1lPupZHMT4aot1+g69nKLp9a/Y+bDndVpnA/2LsOLZL7Q
Nk2Hv7BVAsmSuxQhwSiApTOIB1qn5GT1WFll8Ej40c/k8d/gAEA4TtiGYDZPgv2M
5FPV1QQRr8jkQerzj4/8zkzrDXSnKe+9gtlJCtzkNL7WJsKIVk55KdF7TXtZhdUH
CX86zh4j8ao17rPGfAQ0ejtk0Ib1YSyFzzfxwTmgakHhoFZhJz7a+9c3EAJdI9In
Xrs6mgE2W4Nx1VSRIaCAPUhUdp6hIx8XvsOeMra6QsOa5MWFP/amP3xIgW0DojtB
z6OdidUVOb/Wc5AMLxUG20RX7dFwI9ClAb2Ycks2HNBsI/EbgxUyYOK4tonoIgeM
J6nBGwKvCXnx4A79tlfIMPWmW9BV13GDQjfw34EzZM887Jrl+vuyb1Lg1OuuOJG7
HYnm21frIWCfmIAuJFueQsa9rhuT7SBnGWt3wfCEjkIWoGragyNjPJWNdm2lBtqD
vy/vYNnJWSLivQfwl1XcEDj+A0TBz7QgC9gu8G719Dc0gHN1eZAdhZxzWKDXZkXb
qQkVBAFTDBRKfqZVtwPqktMVWcm65RitoWbCqRe8e+OYfyfBX7KOgHS72EH6UnP+
jThnkZYfzPqBQr7IA1aFL8+fUwqR+QubsxOQuAsbvpAid2Ks2eTeTyuyM017AOu3
5zHL4Scs2S3jUMjbZhrhThL7Ev2PDRa/CbYOBrrDW12qxQV/lAyFNFpsLs0W9qut
6JDfKUqpWgcpYUW0u4tf73+iItODMUzyFh66Cb1VHeqrJl+rfa9zYPFiqx6vlJnb
AJQ39vpbGnW09vxU/avEOvqM4CRSsPU1tyKX/AqDiNr2xCW+MtzLnSUPkmyXvhIS
OO+zIomzkPI4LZrRlTE2nie9IpbTOhdL+Qa3j1m17gzRD5hnA7QudD+sYAYvlLtr
j3Du7aK+rDAZ9PCJLCaGRS2CoZMSSJvwC/NKfVjdgyuJux0W5DfyQy0yARJpJD3N
6Ke14c//MQYjOGaC8NUglA4cJ4k9LhDQFd2Awo7w3zTf/cS/3KfZH/Giqqlb++ty
en3mKSa1vWLVb/BFcT22cOFS6usb95PziuLhEMPJJH7qJMDFIxtyRmuJTT+hVup5
cJcT/6oQ44gEmJALLmIoDYECMhUqa5JRCPw9deboxx6Ni1sP6A1Ghds/Lvul/KoY
KNpP8232fiCu2olPFH0Yr7/BxbWtxS65En8aHZ21xI+TExjnUN6v4ozGwDTFWurn
MAA2X2n2MjbNpRKTXvyKntJjgYF7kXZ5sQDkgSa1Ox3jnoxwPRj+xBCdcAMDShH3
9LLdEVy9de4ZdabtHntS3QPgTY+bKZdo1YUQ6DDzOFtSveVblXqVClqlrx++ScL7
H/NzJ7rWl91sanSgxmJhFEn9+q6fhxJIra9/PT/f5r1LlZEBwIDpvV8LEYdoO2+k
AGTtXcPAoflVK6dS9lI5h1ZF8ywzwI6no6U/CAZPdQsVAnkU4CXALAihc5shBIcx
C00/0ORAJV9L6m7dHph+Qnw4/CmO3K9fNmgnEqkc1AK6ZoDBxJQvQimjIYuNDlje
v9ZtzfHgkZQgc2Hi6G0Z9Ebz4tzEa4wPU1uFGjLneKeqmUVogpLPLNWxjc0yn650
+3tLzqqrw0oJcBYqBmYm6lw8lHv4bhgjC8bUBEnbS4LH6q30LimwYAWCETz8N/xV
rOdq1Ih7d1QEuIv71vGuT9MBObuOUjYkoufDqOGqkZ+bL3/OHoXTkTua0jhz3tTc
ilMi+n8gxBv+490lU/ipJsoBY4th6nB0PD8H/uvpTWjI9cBQRFk7J8NUmEAPEvHp
KDJr5Ax4EpvmV/NhpdOEaDQzEupharjKu31riUm4qGghCUMRwwwFsuZZfTgUpc0W
FkmMuIbc22j+Y4yNPtzrQp6zGurdmX0MaJ/dSr8/tz2W7w1cXF3kGTwdCGw4LhYs
ZKCrFzAZvWwURoHUHwasiLJFHhX2P04pfzkFDD/xYViaWz6dxWv4lBJxbgizhyl2
bEswRly75zDNFNTY5nvM3c9nStkabQu7VojYWA2s3BydEBV4VMWkPB0DVwznsw+n
9Jj4bEcl8Qnvr61PnMfgXpkNBIJZIdwpy+/9/iBDgJWIXhJXVL1KwcqalAzmK7Mt
YUb8CRdY3L1QP7ColPasDDYB5Yd2yMxHXLcsMCiKRo9XPRNZb8Rnq0jzHyuIXv3r
na2mg1P6ijrHJS2JfzDpdgXKqsUnuoOsPV+RKcfUzBOYcnXqHc+0VurhQuAR7rJF
h/v6sIQ5mEkBgKNDv3YLvQhqzELBGckL0tPOeVc6S1mdF8iNpsImXTlEjk7F4Ykv
cCQc6wwi/cXWWhVwHHccwiXEy3o+Y6rT+4NV++EixJkNx1f/MEwn4Inw95dfq9VR
KJqPTTu8m2JQgpu64i4I/WoZccs4HNd68e5ZNfWu9r1QFuqNytW4MAIvWLuzo7nM
iMtTmxo6Xl/iQb8Mx8hcHMNiCmT3aRxRZrMfqITUiBMYGzmxLo22Otxr3pmF9KIN
k1uYTeHRfMKr5Yp0w3uLWODV27osl9ZQLIY2ilV1eZJDfeVwv2FYE5mUGxlViRuC
hmmOOoXkYTWIJnUlsS1sj4lFhi2kPjFyhRpfKZIgb4LruLmXu91LfEqrcDeJkbwg
NXpryYmSTGC4eyXxqSBtV7YdF9Sk8r/ZXnspWdaLAf3HYkzld+xBq6+d0X35r1nO
FtuxLqmopJefkpSinD2NIgcJs8Lw541Fvfwq3mUpC7OJN1SZS/QUa2Ku8FiHo+cJ
QcKddipqBOEPYFXj6TQixWuAsu75u5ZyGA1ajx+uzs0qGts7U78yFwGJB0rVTOzp
V5MAbxK+EJma08074XeM96HJWfMEGM/EiACPSE3Kd/dLtYN3LaVm6Y8d4LFwggRy
B56glksxpKXtWdCXvw8kQVMX9x9aNLe4TIbuxr5LCUe+6GoqmpVgIvLnB98m7pZ1
NngnRjVgYZP7TtvmvSfWQTTYP6K3rkSLL/glrWbxk8Exs934o+N1NQDuufuqf7GY
wwEEh3Tsn5QHltjdF6h4Z9HLP50U+HsysAwX22bTvcZHz36cWaAusMZWqWO/LCcK
6EusIaXafGb7tE1a6WxAnacm8YUtuHHLARl8suvUeJiuDXr9oH6cNsB4asRRbdSv
CDh/CXAMpylRAfT44aRrXYR1GztXwettK+9FCF0C1zzg5U5DaPQIdYOr66nU4b+5
QWRVBUBaCEHI7oUYkbjn3ATk5RtsZQOmb0SPDtmWYrjKAB/k3TnNRqsFoJQSRd8y
YCrp/38MgkQhFRHAKm2wKitqzGIBmjycFjkMzqOLS9UEZ5mHoalYQWTyibejCyXb
IHxPSoKRqXz+j9zDQJC+7r7g/D8L0xfzZuzryOSftdHM3NAo7Wpy/+OBrvyYLMXm
i2OyWWXTP8Tc28DdDafbnbCr1NyfcZ+Koq886gIJgyvuNSS1Js4fz9JxNo7lMeaC
KhzVnzdeyxKpf/3AsrD9QtQ2OwAoqJVSwHOX6M49rpIAk1B77hfSLZYLDO/v9WK1
TcAwnOD52JlMsx5+VeWU3NhkZ1GfM1XpPhp6CqJzsVBe4YFupAgJullGOlbMt7XG
Ty0hypjbZXWQqxD9vdzJZ/PrRU7YXUEKd7x6pg4CizsPsZ59WHRzREstiWb87xX/
UaJ61NNjB7teNtX/2U16ZFC1sRGbL7KYj0GvVfeu1UUzkkoilhklAVLwe/Niq5bN
m8610IRrocoURuH1jP5RF8z3SI3fZyxLyVXGRLJyMxMg/+z1pvzeOuIRmRx8yucr
jNdCVQ+cyPFqS/iXTUDlovIImMOmolC6YGjW+8bPEtMCcLK7YZwqO9+F+5DpwDuM
ozWhbvvsWXM6uEVFxp/CvBK2wxl9XZjT7YE1GXmaPvTG/z8/NC077UhgV/7tH87o
oLk70Y80eHl3YY6vsuYmq55aVpsifqp2aDx72KjTofsYvOlwjvcIwDuwdGc9HHdY
GxnS6+/qGh8eReYyGlVvqz5AGeEkjiEVFszyyGAqvKdrTnKmswxTxm+ETvY7446c
ymmYe14At5sojrVeOiy3VceRrGBUeqffWRKL84gfSTwD7g0S8H5POShbFMApjFiX
f9jzkp3o0J6kFGmnIKaWFskcRQPh+KPMYJAnzn14B7yEENJh1jVmV6ynwaa7mdV1
gw0sE5UJDD0QDIy1UUbo/qf8hGvG7Tfij5tr8zp+EId3OL0w0N9hbt2w6cRvhyfM
4b3O/9n7tXeJlRoOiki/vb1WXFjOmPTk0kJUE8NjgDhikP1IpnEM03W4QRHXWdTT
mOSofz5kuU82ebPeyD8eviyHmjFv788Ejnm28HwUcYawS/a/X3vuuP/ufqP/Z+4v
AImxpKC/i0TYVbI+HcKph6atxIo66RXPlHknoIj/h/HlRxAqnwnYZANmel5ONWCa
2+mCRA56vC3StDZ4Vtev5TaBM9LSJiXRnikGv3nhjpumNvBfNieLeAGk6hzD+mRM
3x7O7u881viCDQixFC2wJINEZhcBw9tjpjjFIY9Vxnkjt6xEqhVJbo+dWzOH/YoL
Lk8F3/tZ90fTxojAXYM8BPnNfg63qI4TkYJkUMw+G8grLaTED27CtQ3fU/UA3nnc
vMRCJxvUo17mNxHia8YZ0PWODNjuLPeYVIkN+GiEbN2Y9+8dv1TQ6sxeOy+d80E+
D2Eamg7CRkBIjZc/dLcVplpV97GyzGGetelmOAG5b4m2DVNCqpTd/tHq7MaMvcQN
7uv6OrFR6x/2mNlI6ZwPBEDdkCi7AniDxbbJUwQxpGluXgZqN7uzX7wo4HNyqIs9
oOZqh2wBmiASdzNjv7TwIYF6Dwj3DboKeLeKCYd4H7zitNpTfM1TYtJbT0v6r6ED
W3BtwqzIrlok0dDjN35I2HgmVvGixfHT+eYK3cU81frvdPO0DDasfFNWLH/akgmb
7a8FvEjhDVD/JzCQ7F+RGcV99it6wQIEATrdm2txQ40iMtlPiDWYTGx/bITnG6Ks
AGYiAGVUyXQcQIlo6VtZMI6o7Ph14mbu3Kytjhz8bnS/ieOA69m9y4XRpOLAd3wp
mNhU5RkKGVo72HSHSw6u2rPVpEbRqqMe6oqRSXQvhC+d2PB3dkls7ki8eo8AdCPW
17s6/fhy6I5jRqaTTAK4kOWExORYch4qoInKweFNP4MvfxXTajHK1YIquJiAFDMt
WpaYM75aqsqVc9367D+kD9JDGyiCUe0QUuW07taQdZ1bpGC/3RKOwPUAR1kMhQ0A
4r7ec771KUrNB8MHZ0Fgd2zIsytnxBwACNV7dkRV7Sa7dIgOMgtEDdcdVqng8wSr
YBT+F6nqCoybOEG4ixGyzj6SCsCZjNdhM8+63zhbuZIioHu4DwR3YPa1PDGjMY90
bnHhxHj2E+EvNrrX+UzTzwAFfYVH6oB824h713P0RohdHgAI2ZguQidE13d47xeX
9hu1+htjKiYZwN6v+CkL2ixBps6S21pGmF72xCdkYQEBVOp4W17D/rRHYb1lqVZ7
HDnp9GL2WFLdXzEJsduoHmuaN7HTxo7N9XEezkxv4uUkaovPnTo+tCGkstWtTgZp
1e+6EgSRINIQdtgr2JyVhMGBgpBWLme9mg6LuK9ngR4LDXvN1aQt9KuOs6D39qhL
YAuw6jFCx2pvpBwti6h4y9F0lDJkrI3vEQ0C7RmHStgw7ONcZKHT4hnp70Fx/OT+
k/TwILSv96F1xOT2ZjWe+biHvY/9cu0d1m07jnRxn9RIakCXXZifdplbevJ/En1P
hrv2ymJdTXWWuj9PYltPe16RyVgLNvF0F8EJEhryuKJtprsJED5m/DF5ujPlJuXW
PN24pHYgD1gkKCtEX1RlBqHZY0O1fTVl1Ee5ra1X+vqPSp1YT6RbVHJdC51vEods
xM53/7yzkz6eGxB8qHQoGF735ebVd3n6CwvgVDe9ltjhkG372zOmyvEwgwsqWKxi
L4ujpdcWEeb2CZJ11RQcyEfx4oBNgQdyMtKB0fFUdzOdv70OqfLoqn4rdgqm4+1g
RbC9tuaEPqMmkSaY56bbTqo1ESSGM9TFmLtui1AQenljQ5/NkrXYV34JEcQS3SiC
aAmq2LHpgOWhmD7H2JaNoBLdlM1/mbGF7CHQpk4qRJRPoBBrtqyV/oRQxnUZf2z6
kNfSNpiMeptGsk8GsAjWbQ/VVueZEvkst9LuAH0pu0sOC+fQLzQQQOK0mq62efMw
WvbWlHwes+MioWCOGD6fjTd2VLWqwLLJ/9197aD6nqr7vtNm7cnLj9WwQ55UO/fP
9ycyI5vz1Ty7WMCXr3obJdANMRTcE9/pCROY+9uBS+XSaL+J0d2mVq7d8a6uJOqF
mtwH7Bk8WCWF3VhQXqMmWdi64ChHCw/E6OdkIx0MFUD0m7Kf5maQuby0Do8m65NL
4Iu36kTShxMoB2Kime3RlklDBdVpgC79qxsTMXb3BlMX86v4jGyKrkHd7JZiTVlM
9croDpAyemVoe4NpWj/Q97ofQk6+A4g1r+L25YArtDSia+uS6xoTytGLgQ3bbWTc
53Mdvqv4mWHR/LrJETEhnsG1BZR+JH8ObG6kXOjaNog4m8VwjpeymoQEnBVADZ6m
j3XLno0tchlCnoOgwj7Jy5apZ8T0rEhJTkWXopRdIT4m2xbA21fx06B1HH6s55VB
DDPrtuSfTEv05X1v/BK2KK0qyT3Bn7xVGp20pI117kQ8ews8Hvftc6fHpiZSY+es
I1vKguEeY7x7j1cx3Y8LoQ/TmSVcwvBQJm2R2rexLVriPPCIHpP+cbhmCXYRjN/i
Ln/kPZhYdiYv2CC6KRifbc+ltl89uAIaS2twyCyF2oeqdrVqWwMY2OC4xP3oGRrg
Ta5LWy00uIJ6KyF63LTe+P+00wg4NWh0WIul7CMsOWHw57ufC+Fr6iWUbgREcPMm
WqkPYX7urGDx/WTi2uZH08lhaFaFiTYdswBZ9c4u/r4rIbhb0N8BZkla+cKEYsqM
mq64duHSPyZ8b1wrTrLTJBZqV35svN5QOTID3rrw7FWEAAfawJK0nGwUdCpRoHfe
GKu1PqEtbbGQ9uKhp5WAb/HT7VcQ/z9huAitSc6iiH6MuiLGRdRrN9xHm8OAjbcp
xvj1+2/0RM6F6puWNDMLoDc2yOUKUZFPxU+3vuLEzbkaZmADLNh6Q+Xr6cVgOpHq
kcTqLH9ddy34FcXiurcbEjBofoQ+lLu90rmyvZ+7fQ2TPfy0KMGlQ+NEcldrfoUo
JXFzhfubREkx+rLwG5HVwdxfpQdwybH2Ax+2ZVSATuchcYeigvGT6mAyQq85z+v+
9MKUHp2L0GzzJ9ZOpq1CLg2FzQapv5nNb6dfODdQvTE+gW3tyAEHzbMejyhhMwA+
/M/AQI/sYbsAPcLAHLjIpdG97C8sFYvULVw7EQIxe+MGc3A6H7N5Ptpfl88uqSsX
twbwfsY5nhs0rVpuZDMfBkW9ocrEV8Qnfw/N3XgsFasOPN/tXh310gV69PzXJXY4
RuvfbGRYqYm3SLHMPCBV7cO2Ml125SUolA6+AACZ+j7/TBzxCF+kOJ4K5BOG+YLh
j1M/vc9cOWs1m0ey06UP/yYryPodeYc2BYHc6ekvCtVmXckhEdY2zdRiv7AX5VvE
gKGlZUuAwb5svkeVnvD+skP2Pt20fPLPpL7bquzyeBP/qEgbCWeTAtouNyoxpeQA
9az2hGpdv/sKRuxUT3PQBXdzu+xnh2TBw0EKAD5KCi6O+CZtVBaUKcscX42pcE41
rTBNPFSjJExOBK8rjv6Zxjfchml9ccrIK3Q7zmnltoFjOangU50WDrBbq4A79WCv
EVKKdUphwahAOSoaSPoK0UYRjhV1+7WJrDMINNfBvol7NFCD44+eFBUmGVxjC0ea
2nRH1B0JMcYlgjQLOx1rLthoaysyG18P9wtovNqoFUnsMK1/RsFjWw31one37H2Q
aYGuxgzyvzD/FVKws69vj6U1IEwsLPw4TPfpMksNRXhKokfrWB5dBAkK3LCi7zMz
8nUT6nH3EXjRtIiVFnxOyI2t0UPTVwB+ZSWHX9TJaDKqPGP3Y+la+LyLBcwbbii4
if2fY60264uXNereWVhOza6Nc3t0HKM4o23lx9ASP76nQY4laXJTBZNOZz+y3Fqy
vq2hsXUi0QS5pfMQjAZRWctlfpJW8anX7q8VXTMfk0Pv+lw9ym/K6UY8VXcov4hi
KyH7fd1H7TOXr1gswGI6H1VxS0po1pEzd9k0QL4+T8bmZlLdSZWT347ndyiHMyd2
kLov/aPwwE20oJK2z+PucX3Bbzo1VW7fS5LgZlfpHWDM9GmyUAFi2IS/BHO4gXNK
Qpj2i3SrUl3Cc05grq+4A3x3U4kK7FS6y4/N35krqcVl+vXi6wFel7iZ9hWEBQM+
UxRfvxUruiWbuHwQf43yJE3tefzDyonX0yy68EedijS2T4d9xLLLKucSddvYl9aB
gd8H8UPdLh0XCInIp9uCihXsesM6bfS7AcYQHqCcejKWjTijIXSPFhk5ivnWWIsF
VUJvETCKxs+ItZykIIKCUXbE6xqZh4yaD8yr80aJwT7uiChOsDMjy2H+oTSVoaKV
0pnEWVSBwc+iDk9wNs8RgXVrBXoI9/U8B2EtiHj9BYTlsgiCTRRm5MVdehsQW5UK
MZ9aet0uOTrOwD6hnQ3dmEX8C7D9vL8V8PL3rW8R83vMywDLwK9N0okBW6U0DKgL
C2sPuf/6HnaQSICaVs0Ez8pTC/Fxr2eVlkpRlZVVUnmB3wyiqxHuam9qokvLiXRC
k8gVP8pLmI8pN0dWKNM5FQGmszuVl01AHm+Z4I1dI9YwGAH2gTUD6K6ZzaFt89wL
2Rtkcq7wLdcrR+HaODHuf6QJFgGh9gF7QWagjFM26pCw7xArfcBkMCrdSfXHxig7
QRIBj2xbvaalYOaEZW0vRxAD9M9F8XhYfJPDUZODVzP2OXsKXQrwUXflN5yWaPdw
itT99GxC1PJQLXZGv1mYtbNNi2IYJQOOPRp9yR0cQqoESWAt28dHTpiZ8jGy+X/m
hpYD/e4O9tqhzQRGmepcIDaI8FmgrOkWSKJq3xZW9RbVUtdEM69p3LaZU5m2Assx
SrksvTJmdqlnWZprHs58455B/X9uL7Ka6HdhPuu1X9qkWzlFVYUetUTxKci+gnWX
C1BnWQAUId6SaLkU+QRl142CEC9WmI3FxKO7ULh1ZECuNaifTrjyvy0ken5PmiOT
xv7Js/ecM9sL5855IH/2HqEZP5aNpj7K3AQXA4zDxADLJGI3NJVl78gTIedoEVQT
sF1AIlJtVcTvBXaPPxyZy+W363PnNFVQqRYDmd3KZygbtYdeItsxPBoj8pjh+TBc
ZBSgje12HfcFTaM2/0tDqnRKDWuccqCddVod1WvreceGh7JpkoQ5PpGstP3hQHxa
WKz/wuKHA91DC+ULgAf6pJOVHtQVSeNJH7N74G4LlvToys4jAm0//HDWRmoMGuyL
ZtSo+EuDZgZgVOoUJ7dbF6KDnZcyLFZ8B5mPssLfy+beDPGKll7M0kx/YqIyaQ9O
44ftVgJPxvJON/jwz/FJbxnprNUTNN+vWKkP5qUceBbpPyrD9VQXyHVbMynaHNf/
Hx0zyK4yeJtAEk3LCXKcYxzvMAKFEcQUBgTE6S9xUmo88J9pRV1s20LtIQkv+vDj
DVvbjhHrqD07173KwZ3m1lNCM9o1Gbcf+bH6Lbf1Q1khsCQlW/OK8rvzj8z/Ilus
xXpuZw7tsHKYXq9/OMeUBFADxrL6pHwvv9DIm/blZNxu9RO+vWs5L1jckBlkLZjj
twXSeR2KjmqxuY8XdNwWQjHKHRj9Wi+AhYBQre1cn69p5a1L3kJA26Z5wIlrJmbI
mHNlxiE/aVXwdKMqsD62eEgwpr93GAZ6bB9PizA80JkKgUCDFvPnNNj9ymiSzvg/
a0PUKH93a3RRxYkTXUkB/4+eMUDghRQdlvtWlt8tKgeg90jHVxNL4gb8YN1pjMtG
PgSbbhaJyhHWzQIC4CwrOTS6bO57N498scZDNVp+xB6CGCTDrl+UPVp0jDi2MDzM
gmYEL+TTx43gaoaiuIqSD9MMIPgGHA/QeM5WdTUr9y6zRGyuvh7CF2zJCKf6cCI7
SkanFsfkpPsRWwa7WkCU+Jr36O2PHh6/Q6oKq1x17qIsToAyjqXgm1P6NDKdI944
ptFDOrijYBYo/cFA2th+D8qC1y4I+dNDlgg46Jf7L3x1fDK3RdRvkSwZqvxAEUgr
I3MRXCXnVrAs4oLoshr5IEqq3duETPTixDBZsnYs4Roxgr7nVRzU/CFqJkU/ovus
4kys1VMZP0RYCrmLEbAfymAU+LaDuTTNi9j6rz6u9qYZr2/c0LW2Um0g3dPUlbr+
eNoumC+tlCf5lc9AsaP3hajGys4ACAI+nr8z36XyRdwMtDMoYToz4Hkkqqmf092A
30o3QLHILXnK8tjdN8XGdifpRANgd0zdDASWYRC/z+qXc0hxH/i5B01CjYn5gqol
kTxL+vEF7yfdpTxpVrGN8cABthWnLAquu8DoPKUQxiKzPX/r4rQRoASTrOVEe42L
a/ZolbxoAmvu2j4+2t5iWJAg7IYFbgIHA5rC7s83pMlgMLIcw4W38aDVQZepIA6E
QGU08n+OtBkbwOiX/0JsQvojvxim+XM1qmFBMmLguhusRKJW09xCKwnNSa2P84BT
7j1mtnYEheF8fGdJ4uYPqZZoVs1JtOEBNE291xBoioaMqbDnQL3qXWBie1vJpYUO
SnCrGHU4N4YyFPAnyeGNiiuhJ0rlpAA4WEQqrxETsyvdi0ewyTsmHrZvEtm9LFMH
oUKY726mLFGyimje4ZadqSqMlT3JmiVD4GrhraAeSbgqJI8OCRpuWwzMG/ceQCVC
+g5ZSpQX00l4UjMdamvlo0od2xfwZ82RsM0ABoHVvu75TqyPQ3+sdAi7kJeGgerQ
DRLyT8qjO6aYKKZSYY4+xiXwotoc767e7nNvRqWxL//zuvV4WjsYVs1XnIaZmyWZ
G95cXNROb/vFDNuaXd0uBh2HxB9cNMePV9plt5DdaVhjxlIrIbCNuOT50UApMlbM
evm6sYFr5giod0+YPewJYZjSJ2OJdQsWBOmxwNLoUhiAaLrUs259ZgHDwFLQnEua
mI5AhGno8wp1Y00bFnxcSvRAM6bbaQYak1TAahyxHsp/2zwdI6lsWCSIre912Jyc
ltX95PZm3UlHIjaeLhL0UTOb84GVqaZXnlECiz3sPwUqeZGH29EHtn/9gSibBC9m
vzPTLWWHgMRyRB+DaRGWWG2mY1aWsGyRr6xeB+1nxEbHYPDb0au7IVKX7EGUCt3n
SOjatEbhOM3vM96A6QYd5VkdPnp7rHXlDJqdRlQmB5SZCSZ3FZim30sR5Cb052+9
tCJdC5B4yjFoy2/0nM+wYmnRqFFWsbPtxne5DWquv1GxbQqBCdkoVmPJxG7EOP7w
gVPMJ8rGEiA/4/DkRh9scRJNf37IntF5COIj/pXM4hhwv1GQhyCcpsiR/P5elOIX
2/5YJ37zyLnGg+tEzuN+eptKGb7fcirkX/bNyFND80D7msxJDX5iJePREsvXnr0l
iM6y4nIxFxrHUvC3Uq1Chc4dSxS9nqeeg2Pve5aKgD5JVehFBHeGteOwWOkZ36Wc
JxvrnSn0rLHRphmBxpw6tD+bNQIrrJdcUIIxUwwuErmxhJfvSe49tVJktfDpvp+m
SfiGjf3IC+KIT8EihbAXbe4r4sNbVHYjrTuLi3E61W2NTWV2jynUY3K6aVS/O6wf
gsmxkCTSL048UupDTmrsx8IimYIND9+WmUZ2kHqGqSRo8oXMB1Cn2oia7GZcW3oT
LgSUhqCYbWMK7HDcH/VfS7vF3pDhxDTpo+EOJldN6D19OC7KA3X0F3bfuFO23SEn
D2MHfFxZqAfr1ONP8Zva8sTkW9IcXGQl3qAF8BAtlJJWWPCnBltcG8ml698K8nza
pVqJSF5cbLblmB2Y2hFRBrvbRiPwzX166u14t/6C1IN9+vkXVoNBHAEQW2FVt66O
qhisfRMb6FwVZmu3/CEbhbRuvcSaOzvNuH1N23ONHAsY7VkqD/SqB3OQXIa2MuQJ
id7gVM1cx0rufk4ZcTrAYmuH0ZLHhTn4O3Nh4r8Qg+77cramiYifzyfT78Mec/Sy
oeyriZJZpPuyWXwJ+IkniuIZhl0t6vP7lj7hyl3XqmxVDhps5fljC2mz1lSgKZuM
FXI/PuCdxzyvnvVf2laMot9Bq8U7ofssdXaI6LnRq+N2z0b37qelluK7VfyFLEuz
/P1R82JTcsuah13JUWXihyu1KNWfnI0v0dXRQ51vHYeuWRf7dKiMDob6oxSCgJYf
H4OFNAIOH5gv/3cdONJDG/D8qBVR3mFx8Gnyz1EWs2JmmY+RkJyJ1FbmDUxoPiOu
dVd1iQLd7CeC5GasPh9PU3z7Cn1H0LJtoLlmU8VhZVt/VjTeG3jlftMrousFzdb9
scMKbIjMDiJqwAc5IBx68YrSgEyitlGInFSfc2UO9EKI9L1Dt/PuScEltuTugrcw
OpjAOLkCunlPRG3sSfuIYIG0FbSkenMSfEhwLqRig9XsYsFXPRGzwTRliykgYG+K
tRaLsjtFv31A789MLnbwcX0BZ4mgFSKglXtgoiJsW3MyNdKNjAp3OubQ5bMr1Mow
PkbBkbiPIaXqmgS3fF1LaFKxvdO6XTJQp+VYA+2h7M6VgPVU8pbH6eCXRSf4nKzl
oP4vxGfOc806jWVwaMRE/6nWrED1CIKYQNtA9n71RnKxDJ32RQcFWH4pHa4sgXBC
4EdtHzN55Z5vC4b2boIZ0IKkeEZFAvp0n2TyZn5nVVj5/ijrXOd+R/4wb12naLqP
JRkts2grd3qOzpr/lRAvGnMcptU1BmkqrXejIkPWnAAMiCdb7Mg1RKkBPinjF0G2
XQiwtFw36t7w9BHOwLTEDS8lxcnNKV+4j8FG0USFWZ5oZlkB7kvSSoCkFcxkea/9
mORW6zyXLdmftk6Y3X5HQvKyUPJnBJ2GfAJMRx1D+MLATbQosknDTTzAxHKZb4VT
oGBp9YpzZtN5hdZbsWIqDTOAiwPim8ksZH5qgBzylOFP+PV4DXRIQqIQXYdzHnyf
E8Q2kQvO/3KKn/mGZNkSlfY3PKanwKKfHxrS1PKb/v+4eP/fvJdBGk6AfVkTJt3y
UekOQM61HztdcLwoad7DV6LOcTIv6S93WShcMbpZmZOtsRJUYGHOLoLIF+FTNaHn
vvwNlvLDJY5UcdPZmgHZGv/WaHDugd++3rFJs29WqEFYpEBGBTHhWjvPtInfp4bt
XMRd6XHy9NHIBUCyrnnWBrJXaQC7ILk4nCbt9QrHY92m2aJCs2/7YS8K7tqDSAmw
4g8V2F2ri5cjE9y47fEoRZg6tmQl4JXYYYdjYYtf0IHibBkxBya+ciFfQO6GNg75
J+h0TpPaWKreVSegwCclx/cfBQ9SevcuGRFXVmS70lroG8fGrluKvuu2JvZrV4fD
o2mQvBSGCReHK02+ex7h7sJyOZiSM6LW0UBbl+WEVkswCtDEOJAtoh1lIIWJDsx4
rmaJjYMTFxEDrMWSKVbWJL/ttGf7rg5kYfLolDLo08/cO/tVVdl2bAHZWLOTherN
Jnhm+ddvqJX6U7IZRQHmolYgPVaVePMcz6n7aSe8xmbF1500f4pjI1WUms4i0wDN
w8s0h6kmZ6jaRaEGVjfap5S53JYs7h2ERbTEstXC7jKSLt8R+w84hGo8P0Azd5HG
ijEqeQX0mBLvB0EhNmIJJCHaPEhT4LSultyOmzYIXPZnfktjAOzladvBwIdAUSLJ
kolA1azXqyDnkxJRxHUAk/QLtn3xYQLmkd1uDLZVaX3pGSrGrs+95GfLe397yVN2
atksyxc2cjyZx6bR7wJ6AgGs6EbF16IYlXWdSG+jvAJbmcM8bhpwuGA/hQVPECrR
Ewib/uAaomTYLc26SJ8rp17fJwnKKEAD5nywGgDPY+fBz/7ccTARME+pkHLd7OxU
pQexHRguS6SM82HFd7Tv9W9Zs2gU4KqVMga/623jnw/b5PN5Cka79NPN9wDVeJI1
G5dxvtLLqb4KX5wrCNgh+DafpiQesw8E0q4aKshYXxCWzBMHphC9LjLRxsFiw06p
ngCbk6ElTK9gn3MGic2oft0jBVUi0Df4/eNA+3bM90r0fMRLxKW4hagAq7FPjS04
ZGRliFmHse/rxIm/gRobrMYW1EVF8yEhuDe89K88KvtNLe9hcxNv0RXPC/nwlMHW
Y0TcdQkzY/7/EZHL1dOhOe6BhejQz+hNRDxkR28/hfQy5GYesMynGjjTyYFXEkar
Mi+Qepa4UwcKvj/pd3QojdE7WtFkxtfq9s2xzztCZxGr/B072tv9xqbbF6JvAsWc
XtdCH8XpFat5jZMV9JpcNI3QT8kZ5/D9mlw21VUPO9lzqRoGQLsBAo1mTkW2F+cP
OQLPrD0XJ/ATrtdFNlSC3uuoCQUSJhgihhzWkqypet4Jw+t2xglt9Kh+TZzGNvsp
eTnrp63STzEa4KIf3fCEk+VxJVuwkyKCHtUuEqzhmQklk5ODyC/syCa9gjsY4TJ3
IHaQUZM6dz13/42MxKsoduC23+4zbBW9yxKPyfwp3fpAlmRvuAoNTZ0cnBvsFIMH
HWKQi159EXYnyOaalXzQo9IauiDCweXHMiD8PeQMGNlB9IJp3E6wjj51m6Nqpaha
upHV33f8KkfbrokLItfj12AvMDhKCiqPIcZBd9KorZNDOsk0uFCd8Cx3S56uP+Kb
gZFFf6pa7AbrAN9+HnKXM+m753sFAWVLdmlxYEU72WTK3iI+Zui+wxoVhdUTY1dh
H0u4/b+4/99taS2oMy80KGp6FoiZmeKie+TFgS99EPrTaBQeDKA3gx5WcMKtGDIK
0calI3TLQKpdVkKsk2uIO2UEZ+7WDDNSRXpmKRtvUgOP2Y7pEi9HO2oIfwBBnOD7
7LdqYBGFDUyjo+4cutuocWanKXviHQfR+ZBgFRktd10x9TdqJsW5l9bFPj2jhNKL
erJFNSFoBJ+Kwr9yGbVxWiabMaSALwUZ0ygrsoHtcXxCG7sxaSL32UsLhADmcFbL
ZH5S4zi57kKKG2h8B7N0tC8QQZ6oEXkDv/ii3ueRoFKGyKpHA6xCQSX0krgGzjcH
2YQREKakiHlIy3lRFgPsJTMBRHHAEhSpLhJMvZSfpwB++e8gay0lClhfzlSjwAzf
+vQ0pTr8aldV6KxFnz8OLwAkLo0uxTk5fOurKRjhoFsGA6EaP0dxpNAJrObjpdeu
txozyj93J3+qw/dCKuNUItFnN+wKY9Bvf5WZc4ndnflOSgYWk/LFLjYFK9Znd7vZ
h0NWlWlqLQBTyZHYIOePda0GIoiA/M0aEMX/bAXL5rzsJxMvz4dvaPNp6TcgVD2Z
slh8Ov8XrPXj0sEk82lmhg==
`pragma protect end_protected

`endif // `ifndef _VF_AXI_SLV_HNDLR_SV_


