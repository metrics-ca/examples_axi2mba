//----------------------------------------------------------------------
/**
 * @file vsl_am.sv
 * @brief Defines VSL Allocation Manager class.
 *
 * This file contains the following VSL Allocation Manager related classes.
 * - VSL Allocation Manager class
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_AM_SV_
`define _VSL_AM_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
myH1prNNl2MniRRR9snHn2N61DWPbxTFLGUdO1W1ytEmCGaZ71F9yqRahrLih5P0
tE0ihXkLQ5JtA7IlNEoWP2nnm4nzCsLkOcsZG1BBWqbq3WYqvBz/0M8dmEACWy6Z
St/6V1pQG9SxjBEVWeBiCq+wv9r9q9Gytqjp5GVFC2g3Rqjig2h+LHh1NSvQ3dPP
8/cywCJ4+7xztIeS4s6vj/Ygh6wtYhTfFlx1lQF2aBD+4lg/y6GVsXC+uqvlxuM7
dXTpQKC9PORoLIDJfqYw0syTjniI/hievwttStfB/Otp6VkW+6spnHCkFGojyk2u
ScaZ6f1oX1Hf/N1YdGiD+w==
`pragma protect data_block
1p3qLUtUyrbIB0CVAKiXdrFZDqbz+XkULP/+wXHzn8GC13ohAlGu6Ca5JNvSq26+
T0NOS4sn8aoRO5DoMZy0KR9lcQuu9qBRhYLNglvpoPckcqstXlefJrLcOYT8eZAe
UahPrDVYEIGBFbSGmnPE6WKntN9tg6tD8XsbtGUc8Ok2u5BfgHvExH6e0BwKBIv2
aJevui3Qi9wXDBlTo1pfptBbHcoxLoB1m5KzbTmKou3OEAgAeh9Ub3Jph1nwGix6
CvXJKMWKIKWqvbBqzdtsvT0AUL0hhz8+iixYhQNYZczfIbF8I+sF27LjibtphHdE
Abgr81Mi+m62oz0lD55FW6sP+jfirOz7OPbW/9lIllqF+nOKO5UEuc7zmUME0u5S
9earBtqVFTu/CaljrhKKV4f8O+v5DrYB6ZhlA2qPhDWpmx1Hg7o+nlcl81jufC9o
nBWDAm12WKw3sqhxMKiXOtF8+6IYdy1bqvPlzu6gXAlaxFjwWiOdWjrYswCM9uZM
UN7HvhGZ1BgZ0QA4/QQki+gXYttsVLNItc2HB9L6qMk3Aw5Zn5LHrc84bBgF8Npi
Jjj4D9wF8bvO7UPC32+7AKfZ+5DkW6J1pTXMmop2FWdeniZtnazF4/XIx1lWoTIm
MRyiMWcJNEeaxcabS+YACD1jkC2wklQQd8Vl/uzGcSArkXALfk1JuP2huGh9XmAa
iZeoThPOIjSCiQGlUY3qSs2MYNttEXapbLBDflh5IggqYb/D7Vx1N6hQZ1UR+ILw
bFEJZVKlNAzuZhYXwuFh7xNpW/FCH8h/2j7YTIfeTpE6y57BPSAvg1YYFM55uIrB
NFOdhTh5/GBe4OxpmhsEGiamxzxyWgFcvqn5p8x88mn4/rK6KdwwmZP4i9m0NCcK
wgUr1Ce4/cy/BvOqXGVHzaid9CElgH37xzzXEzC0bgqZZsUgqtxR0ZAFk0jZ/Yek
3G3AQIBzbRptTE0wSoflp1ksFTyjr0J8XSLUgg76AtG2akNC1htvNvUCQnfA4gB1
0wfQwuoT0S3/0Lf7K2LIoOLfZU2w3Q5V17oUrWzVRN4oNkwEXqsq0R8sugjBDXv3
Heoz/ij4DNC4Z8CfA7KB3LdCQy6jz/a4lsdKt9Yl1J5nLatUiQ3vgsacvFNbd8An
P+OTuJkS7H/gEZDa9j/Fnl9zZ8bZPKW4x+h/z5u3lGflcjsciLLc5L4j2z6KGyRs
XGvGsK09y9Ob7JkEeUZEgX2W93/BZZQkpy36i1F7hcMG4ODMxHT5n0yB7+vIydhZ
mguhLz4eaBg2T6m2JpnJd3qHGz25VHbpPr8r5cLe/1sFxmlh9hGbLiUhG2XFRWQO
NVoSCZI4BY68FFQwCCf9TNZFPHvki/VkYpGjAbWbmnSn0WRjSlmYoLlhbQHrfn4m
BTHawjP7xgSE5Vqoe7WnMkpzDv2EkUFubH4VhJXcBWcDJvX2i2Up+TLQGOvFy9SQ
xdpYDQVd1pOzDpzXokXGkcNcnvpMKVSu7iLG+4XmaSWHD11uNv+RAjQcVawH6K+A
SR6WofIAjsJVExwl/zWItODtV7mvPec0Q0HKzUgvn0Xo3bK9wgE2qFD0f7kwHvpc
8GzZDBBMZdnUT7N1oRfICFAbY53iPCogQL509cZ4ADDjWLE5Ov6cBy087RIIQzIm
Dwdgi5HCrnfainhOUSpG7jfprL4lZt/d4WCSHs1aGoItJfc9Jnr/0K3dVcFQWeNB
G/Zl6u03JDvyIG0dtT+903LXaCbpE7jCqzdamyNOnWIgQnc56nv/loHUJYVGtxA8
5GwvH7owEGIjZMd83q4QdgIXgQFBQsXeoSP3MHZ6ZNsQCnoBVERkQwAnStY7Vz5W
rijI2bkFkTUPcHyss7XUEi5I/BO7YYRvKMrdcCXo1XdXeckaNbYzoV9o1AsiK7GW
WS0/kkF6bUVKJhHFi1hSYtfoWaHDygTdnSTdnP4OqJ8K700HBUtG4TYmkYIZObS2
WZVtJKzSwjBzwCiSpNK8YAETZcnZZ9RNtvY/ZOhMNXGgmtl5rKWIwrrDR9Bl17Wy
erHZWTS9io6j+UkDKtldfxIXv7gNjkeDLFt7mWm47O58WpJo37p1q6EesnCImdJ8
u/LFvH/FjwRKcwus5XwbucvAUcyMdVYXE0muIY0JA0DuOKayvXsswe1SS6TB372r
d/kUm7p+wNOcx/+aNIFG4m7a+4/P6RbJhVV+0nFnQ+HOd1Lz9sVCFpeMIBpOqVZk
jkRuqRS10sVvuI7TfEouC1E2OHZCGfw7Bcty6oRbZOcEIuJ2aBw0QSlHI38Nlfbc
ePZwsROWM0g9wxozCo5/0SvJSNkGOb6v1WENz/fa7qsbWeI1vDhmt1vVsT+3EUh4
ab1E6vX8Ui0q2SIHLkrQA+FjVzJUdHrHSIdVHNyQXm1u1ZsHwS2b3YKIomW/EaPA
Wkk/5UkWu9oKO5NMGLwaYQVLoSynANi13OQqR30Nlzs1lw3Ur8ARruLFuMXMAHyj
UetMlrQooCZMdlIR3fGHMPYp0XQnCkZ3WiXw+hkITbxsybi4LDRicCYQrhq1E7qy
h9km5f99YCcHCKcux2N6aXFjh4ZEHX3NSdqOIcBu+Fob2MC7bn3dVVqRTDORfSOM
IxiJA5D6EqsCXMYamswu043lLA7RvixFpKDSHWX2tFalMg41D6Ahy9fal/3XZQr5
yiXQMMABg99thrrHASdR9BSkb3VCH5Zax52f9hyPrGL1DEZ2f4y40EM60DNzfd5z
5W3zOHpMI4yrSXvOAVJavIRtC+FZptHPU4BnHIb6P5fV6VIMpBGfzCgLa93Yasyw
gWMYhafGtlZt7sG3HerhFxlPvwWU+O6rG9+0T46ApGKtgoa/oKo4A6s5oddHhqSI
UmYJGT37g+2TnPXk7JvP/qvdWz5dYIjMyEoxvPdFlfuSpJ+Qg7ErRegrMu/2Ax1e
fqG2NZ8IkOyYojBk0UoK8weHbOKFVjRCy0dCyOzz94NDoPKlphV3hqLYlJcF8srH
4xME5y5wIMZEekc+vExoAYb20IScAToEaek7ABloQzn55xFtjJ8xdoJsyIdyJgBK
JBI/y49d32HDFk+ItT6OSCg7zoD63cPBJesT0jGm+Wf7OQRI0/HBCr9gtcWwYf8n
fCD2jAxhjEb9RtMDWwra7YHiU2RQN1LD+sJdw4u5xIhhCqnrRT5v4C4szjyLcoCa
Tm8dDQE2lLWxOxWcLz3jivJ7PHwD3E9gtVeUn8s+PhWkn6qikITD11GEt9xvz4mk
qObTeaeLrnUN94HleArv105+50/nZTsnOPr4wD1SfdU9v/DmJWuh886lYCpwq1B0
r1whdjLyTSVG6RZ3fVKULM8NH5JD5Vf2AD+PS/3GJGeHHt0X4BZeMX2yVnFcQHw2
zXv3GgqHpxhP6ZuTEozBoZmvquQZ0/X75+AcrJC99S8B4jfSgluHgkHIV0B7BZi+
Beu/0pHP9OM0AhQzhby+ydpRliQSYjsTb35EoGocgoHCL+jlqoCnmIXLW//AHzYq
/PxhdlBsfGdTtYzmLd4HF3xCwz7DCHAxSOPQmEB7loCip3/6dHRRmFfm5HlXScm2
+5HbthEr9u0fNjpLPlbQGQekGCnX0UsEhp8HjvGREBFkuoI6shPXRmAbNVXp4RsO
yR+jL3oebcOmDS6vO4j11kjYhV0X0Lp6yqRA5VA6TUDQ82iA+agOvaUlICE+BWNC
1CNJ/x3E4izq62NuLZDsXFS04HHDIeMLwzSHBheDvDnD35Rl/eEDleOkbVyyR90l
7QpNq0ag0MatEuY4mWZGwlT6+KM//wum/B6q9DPwBs3+CiEOeYno1XtZ4CQkaOOh
IGu9C0aVfl/Ue5jKa906kOOaXpGnrYPCoxkUBa+7R3BmIp1UAxpwZ9/SxH5elgqv
HubhJyjinuM3rEVEluT+vDummp5/hliZxqFQbpxtUI3RMY8+1jAxKZT/I1ES1L3B
dz8G6t2dkQ+lpxMNW7lABzEG83Vo+Mhc0abnpzCTcWDVeHwhnuSbndHJVk0TsPOn
dXvvAKEe6trAjUigwv2XO4wYN1c9m3Cbw06PjQdnoAHB689vp143/KLCq7IAdzUA
cW3o8JFFARx0sBcn1P2sBuYDQ0YTEsP/IUCDBRhPJW6ltfrI4V3vvOpk3DhTb3fk
/X0dJms7MzdJS6N9XGAGnXFN8PODFLq4Lqls/yEdGMk2S3g4NjbPB/oXEmHjmb0Z
If3Uy/VBkoTezntfN82F0+acoXB4KhKfu21g+aWtOBcC6vz7RGMe1mTmmeCqzlDm
v7X0b3NQ8SOND9dMunOAJtgL2GbZc+LZ40ZkfZayZ8pb/mFMvDfLVJvSCsn1L4b6
i/V78mrmwGhxsZMarktD6lAtSfw1F3trRviG2RLIIlcteKqG4MUV4QhgQMzXO300
nRzphLimBXL4wYq0jXbkuWtYH90oVxdm1haZUDlXJm03ySk0bEMNKrt+xS7Yt2cT
OIlrN4EdRpiFys+GpmG3ZkHkmqv9t5gJR0rjC7UUHrNo+cTMFt5vLXMclXJ4odjl
xLabjjkN3l0N9vhPeNiJH8dsfOFDJPmSucfL03ndeGPb0txb0zqwxUyI77IEfStK
tEM1jMn1DSqbi+xha5S79u7KshSAFOXbcFo+vsc3lrrSyVbHS1fMsv7UnYHxk2OS
XRIY+R2XXYxgSxGhpx3J8o5MJ/s0FN5AWXte74ChTjsxDbIGy4VCLlX1JnMugkuK
7+5kH/INszqJTedSDNC2OBxzoXkDrBMGBsIrRU+o0aZ7YlkUAvaQQpMIYzBtuRIj
YVLPBN6H8KeTISn9jlZrj8Wg7twSVRhv032hAq1tWwbFnQDbLUw6BHrXN3p4UwD5
SNdOQ2Tv3T72HgtmKNKpZSZqIckzyKPq+4qgKjHcBDlvlK5lvLgUMg6miq3pqAKX
xbG1oB72EfTvH4PAPgByTtU0eXE1qq/RnUyKD3t76iwT96hPBUhmS9CXvTY+47zn
JyYlv12w+pdIOPSKVpME+zW5RdHen3tTTDnTJ5zrUcByaqNAnhAfax64Yc3aCQuW
VGgSCEnaR7EUrihUuql5RU2IJ1TdXqfSw6vaj/x1WsRyYIF0GmQtswW4/A9P47oV
to0ud5fjiaLG9VM2/Gv1HJTUbs3OA3AChi3Ucm5WQWmGSRWz0GuP4+TwFj7B2woY
KLsBwg2edZIBxCkQs/fbd3J7sTTbuF6GPbE6wo8zcTRqGlrWzB9XxhnLzHZ+Ovy0
W+aXdjYWSGhft7ve2g+f4OjMM/7IqbZX9S/SMiRLFShXBcPjlMUK8QOIHRqYtpXm
bErK/Pu9TJ1rtVsMYcA6zW9dxwntCGsiuMZ9XaxdJReqfafCTXMpJRR9LeVhWnWX
/afRUtEqcSQKnEKev4RtmVxWezioJsZfckshI8P62QXJ5wiNFlDcQxF1qv6QijPY
8MTyaoJkzhyiho2BJzm8X8hUfbEsFPQJvAI7+mX6FRxoez+jv87y7AiHAYP8TnZg
VcJUfdkwtPZPqO2CX+xeVrX4sljJKIEzVfZTGZ6vr+knTVaYDqA2numFA2J9fDfv
alRgTxLFmgw7mmCbP/rLNh/w/M/jZIOF413H6ylLT3EIk1d0Ow6Hjd4hZxVHX932
JLJr4SDBcr85dSFwrYrDfh3B6FiAYWbNGOGlSQjiOn4zfAnlrIEqW+Rj2dfdvVJr
GI6k4olA2cQPzTyVMLagUAjc4DyGBPH9QgGpGLbtjM4ZYAetpyM2LmAIV4tDMxVz
kDVaNypC9Sc95VQj1L3nTGpSZfr40eS9CULMIKoHlbw/2ScBkkwIGYHdIBppJ4gw
/RktRtiVhuCHNV5iXCgxZ3xVs3CJKpzG4LGEyobubnCsylcMYf+Q8ne2a7AIWXdD
9Ua7pkhJEbEFYeIHfKt1fNEDkfd84OWzoLGiuctV6NcDY0F5ji39pPvnbtKOk1mj
qOwVrWPNK6u9yOQ2NNS4X9xSvY00DIyOBrMvzA0SbgG4LaFxIJE/gulkTl3urnyz
m5WGvoZLVdupnxgHflvJzItuLEOjiKZcSQGnrWnUwmke1bSWItRcQ980WTNHaAyr
na9wURN7B0vnbtRQXLEb91KjBPOXOHIBoVvSSIGr7SLTj2cIOXbeIUFKygoTnhAv
JvrWXFCvrSf1L/+CU4G7HoaswXRMG7flLU9d8QeeWvx3euO4xLELSrnUyIYgoXOC
Z5J5cDYJP8F49TwFAYzYVfLK6sxMRs6/uJtktRG8iKR5OTmy+18K9Zi+NuJTh+ec
MD72XwFyKKzIOQBn4vHaCA97ReG//Wn2xATunDaDGA9sW30m35gEVIFQ6Bkq3ctG
wTJrTiRfhh5L7+YO5zRfQ772+S4V/zInrMf5Wrk8/GJibTq9xEm3iVamEp9zQh3z
PhWwwfFJ3eWsweR3MumpK7Dh+SsFAlO4ULW4VZhChXmaYQOUpr6ASfKTPF2fJxyw
bT+eyu8nCdBhwNIkUYkyPIZKjAJnqhYZ3FRgiOwfR/C4rpBgfrE+8KsoMsFoHc/N
yWinX/jgU8+1WGEvHNHWEKnXGQNob1GSx5GKhik13+xQOJpBKU4YTvH7PmLqf6ll
VbWRm6yllPyTLblSJYN1HYvSlC2DHr1A7R1v4XtitQia0UoQe8KwLQ3lMwxMqi/T
FkK9vuMyK08cJoQZtmSMRPf5TjV0YIkTqf7QfbYQHxTt2ROlLDYnyA94qvBYh2tF
1BeYUohp3QnNQkCGJbnlGKXPH+YXjdpoQCpCG+eQY+Y88QgDqbSfHEgOnocCKtWJ
D7Hf/rO/sA6b1iW1FuEVPt6L5q09SnLAo0QUZNnEpf/1eKaXUTDIw2vC8uzRJJdg
pseQicqOuFazwFCw1nSVlANxPQ8UO0IX+4REBl6WmHxayg/id3LmmIjZP89nygyS
mFFpPlnwrbZxM2rUs4JNAZcalXBXYhQF45pfZgak2fdKcZUItQb7VRsUYivWuUcw
UhhHXJl4t/li72g/+gVf95ay+bsuZjYuUMC6vSgdeOj6OXNula0896XqlpcuV5lC
aI4UN4bqYPgsz0NxOZZYGPSQrTA9Fz7z0KKywsaPOymYOI9uWrvj3paHy7DR57oa
CoBLlbvGSWcryE0WUj4olKyrKi36ke8nK5rLOl8PUlkVMwCznzae5Fbem/UqmOSe
D3vktg/cYbDNM6fJcyf9i2R6FQT1e2G96sE77A75rAxYOw9oCzgp0afBlb/oREaC
WhCJMxBFp0uG1oLzeEIgUALJMMDmFdyuKUgBfMmbW5dp5sJ7X3F4pJc6Jp9nuo+3
nQHoJHFH5Ja1ZeOdODn6lZMjdMrcIL9z8htdpNZ2JJnN+B1kYxyk1wpeLU42UfuN
ZfMF6vspfV7CDIxi1jvDe15EKW7IaGzq/GLxj4oXbbfLPGG8fg/AGi6rryc0y9ZT
3oYJi0lLc+N0cmf5xysQDRGFl2Kk5jMKMiyeLMOlRo0qf5AqS4+PK1XGnGQCo8hA
RrA0dVGLatgJ9a+tirLUXDllQ2EVhRp6NIv6rmWV/0GvDqrX3GjwzV47fWfGbBzC
G3WzHOTyBcIxvw+K+RiAZkid9MefQHaQciaC504eDVLrClkMb2cuMD70Eytv77oj
M7LrzeVsvTEOewiM2TQHJ4hj8JLgRmD0uISBDmDM9Ypfm0MWdC7BQ2TPvAl3TrhV
4b8BNeSdhWpO2MCFOCU4bUIKPSO2Eys10slMY56gomURTON6TU66nKb6BtfdoaWo
7BIyaQxEA9hKobfuOrVvkkba92hYWv8YaUxJQLo09Fi2fiBUXX+xOyWB1n3rEnjr
1DVxmb0q9lsjLWs/VXO9dHYuqGTFcUJX1v1FNVZjS6ZON9jCS/6N17XlXBv/Bs8Y
mo7wdwxL/e8FXGbX4s3N/jjTAkEbOH2GhmWHSH941xTUmsLc642gkKEJLhzm0taD
TKc0sEGOju9zOuMyjZ5NOBdSrSN9p9jZPIg3Z+jgdsJjgIXq1bVBjpDZReKkAPIO
Jd/hbHklsAPKaJY3x5mxtn/6JgtyxdpRq284f25rijr+4bVofPwNR9LQtj4PMtYK
QCSLRzVHuaNI64nkKbUplpuX+tm1ljRAHpRX2IvYS+W65P0A4VPLqaXH6GyU4Mxp
cPgsQfX0/V8T/Lg8u0ZpWB+QtVhrUQFndzrVZ+HAg2bLqAfbr8GnzF/MRg7GBVQT
AoexNdJYWHxN9KXpdCfcJsTI6OKuXLq8crzFV2/p9N9cyjFE6AVtdHiPu6aGGexj
5PXWKV1RK4wrb307zCkL7n1UiZZROWVfWfo9zt1+XqFVc0d8IAUNHF4gzS2v6Ewh
UoyfRBk0s4TkQjDXaZL5OjcNyrj4ludda0ZYu3IQKfjhwEUcYhcMRBpd/8qOtFZo
W5mQCdPWlDBINpp1cKZveyEYFs3sHFUDoOIzfwpVEDGgjShy8vzu8MjKv7tcczE5
rRrhILWxx80oUzE/xz88MhYrIYDgwBamYtw9oLXayDrDXstjdmiK6hHh/776Dh2C
WC6Iscp4ZdiQypPYn2qTVwO45ZjMRpEoY8rRm9TUr8/ia7EG1JutkW8u9KJRCtNr
SfIyxvinSmBDHXRiEe1IeVixorZiDEKD0VGzl2XOzuTE90plRqUick7SEYknCJY/
KtupAdNfyq4emmQEOaRIeax0Sk7fteLVIqI4aWRm4gzusUKa2w8bTIQdW15lsB3J
1nXiHd88jUxZRRUa0t/N/ppgOnSin0MLXEHj10ceoMqyEdh8QhNGaZmpDsCIxyqA
xZq9A5ahpr0CSW3NPsz+CbWV9ZTMA9b8Vsp0MXat28QZlcPIsX9n083oJ9Uirrr5
ljGfyydsjt0pmLRI/wNt5gp2YKG9LR4Fhthcp+KWxm2pGiI/UVFClIiaYutOSB+d
PNM9H6Hz6QYmXdnvaZxZSdvzlmRealuIY+KfgxqwWRQf46W21ZnaaL5UTVxU1XUC
foC/SJFQreesnN5kN3CLWgAvD5pPe4bcvC94UTgqAzOCbobV+DNKwV2Q4jO1d1Xo
SxpJcjzxO4jF0eE9af9/HXs4lAp6yuZxrSiXu/mERytFjijXcC1p0pYA5kPa4Dlg
kcNDlVmgUMwVgOaPVAnR+wOafRTYQ18dKGxYF2Pzoo20j2xUHq+MsTqXQYfmeI1a
69kGraXFuzZFrbLG+j8Y11Glm0wOL2ok1XBTEAY9wdXwcHM9MyavNxX877yFxqGs
HPUs6Le5tr8mFAXnT+j9iz9Ic5cIcrMigTsQamtJjeIuHhXkVGXKeKyuni8R3Kx0
+chY9EEj9Ir95XFL9eE+dIlkpHpxpTrPRFrqYTdTgeV4sU9s5YXJkL5y1AgizeB2
mdaWV/S/Tl/c8ENWwzcSSKQQ3OXJ6pxRk3FUoGtNbsoBC02p2nia/sPZgdMTrXl0
7PkbnAjj72huTYuj2WQLlyjrF1k+bY8B0vu04lhrqb5R6pk8+d1Hcnm0NXARz7CV
btPjR3qQxENKZGORHAcaFgj6tWz4f5u2VgS/Pqzz8D/ramADQqusNciADT13nmNP
em1fPwp6dtLErfkzpa/MK+Gd7OQiQZbMBgmmF09OshzJEngqqcY4YssnjRoi3IE9
zJc74jgY6j+ncAueuKqupns4U6Fwlxzx52qX39RbpPESP+jZha58kVTidXeJ3YA1
EUhdH4ekqhUJRhsqIUg/Qrcbt76m4XMJe8kvoL07UeCnsiFtx2TYKLqaoK2IFG+4
r/7FfatTKbZE96MBdkdWAMl9z/HWFcmSxxfTktZUkQmFENK9a3f7VoU+vWhujkzI
POlrqolQuJwcNuFMjbr7n7Ls6V+X4ahoo0nNwmSK/eKL4Q/EprhpVVkxMY0GwTdV
XtjJ4u6y5K2KqkwtVbRS1iH3ktvXE8pCfV/7LERW4JNMuBSMh6zASJox0EC8LILI
sEKB4dRNVYT51p9cxdUDRt7k1i5idAUMkLWEnlTkYZEVpB+DJTm9HtxAoEXqRx1j
P4uBb38tkB+iVzGmslyOYSI1n3Y74NHeQK+UGbH/h77R5hMltKt2NJJIdUXTAFX4
ayF9Z874wS7xprNb0wqImuXLdyH72AtIMvNvIkSsagg4T/972KBYH/U5sBih4PR4
DLDtLjNa3XOzQinwyHTZimjbv+Tly8OwwTq2d0/o5C4a17qhR9CtaHCCY/J1Kuos
U3nQAAv9vdkpdzCQEhQH+y3YPsMN04p/QPZQiNSf9IIHLcx6nyKfOf8DB5/l6Qg8
nHhI9WeD4helzQk3pB4UeeFsaF9/1zyBE0y0ihKY+r6cpMnxOx9TZSrxhXjTclCJ
JDaGPUuoQxX4JkMFfUJL4XsDxWVducQGn2HczFM5bNZ7l1LYnWV5EagsgpaqLZzg
1GW8UjAT9vBxIiG7Oy0AzjqwYXCOZ8WmIVaTW/3NY06i5JZIhwW699kFvDyiusuO
i7z7izh5bNET3bw2q/IDJ4aPxdswSmaaKU1lk+sw3AjSQUUV7581ypvkxK6c5PiF
VNulJUVb0d/a542fUs3LnCDGoAcY4Rmw8XBOdD86iWowEKfh8jAoyDzvBxL4jjky
X1XOMfulifdXlThj9Y/gEFyMKOkcn7YLVB1KTrgnigkRaN/MNtXuAvM8KwyEOvoy
17sAO+dkaTIyEj9P+F2n8FvF2bI+4Ow9JnuUYMR6DdtNZCEyuojlkcbASU2QZheG
uk0z/Aeuqgu8Gkf0FcIVRje8ZniD12o9VGmr2uABjbBuYofizRltEtDQWQxLPZ+Z
tpeDau0dGPF0l+Cyw+uF5aBFp6FSMHjnZm88ppc3EckWn9MWGDTf7CKUK8coaUAf
dSsCgKDFc+ib9Zr5rRaVBYgyeTPbYuEMc69Dc/Q/+1rltRLfy8lbtmdFhS3guH0t
MUzSd/xfKnt4KGRh/MzelitLa5/+9jbooRsR3rvQi1V1VvqrWiYiExcd+ZHywNVh
0RpTsX6+xMx6yEAgnEbn7SY9023I7TixRl87YBbHISsdR8QTFkyeDtaJsTXh6EkU
Wf4KNF7+Mw2JQh3/NLpUqCDtDgxqFDrVFhFXEYgG+XaHWVoIgOgFdLr0cIuc/aMP
XN3cQZv+m7OVzsGBAycnrqBY6oeWlJzKsSNGi2I1nwAeYFaorgbxx9VLalSijCnW
FoImchNJ9S1UtmgTXVIBWfbIZxJ1evt2/UHAs+IFGhicwOB2+DIZfaaaQqrr+/yL
Zm800TiObpVPs3BKzeTHDjyUi3ur7IsTcxori4k1rkELhXGXBPZ8LS6CFFO6trx/
qgEie8nGpH1aZYTWd1LO07DV7IcQmAmh6hrxzGEBy750VgVK/Ad+jUA0tTkRCGi+
E5QNW8REX6orE9TrLw91mxGixi2mMtReO5J/QoCeWuEkrDp+0e9HW8l9oHXDyVp/
xJ49pk0RXFAfmux/XYkC321e7Lia/+dRDc3nlREEURYdFAqECIFZKk73ubq9bBhC
oQpSh0eL1urDf4o/l11CrqqM2GtqKnLA2cgGQ1UR1CWXm80icFpg0ZHOQLSMX7Sm
3iRefYzjZIxNx5WIMVGpFa4ay8DF9g4vZNrsfzJpqCTBwZAUVs4paJeq3CXXrF3b
mb0HJI+XmSKu1XJX1TTtrqDwE6rMZbCWQ+uEPGyj4U8q8SfJiYJlEhxlvNqV8K2t
6ueV5dLJWV4C7rfrW6TMPueDZCEFDxMr3XPJU/8yF7xVesG34cXtKkcZAcSiChXv
dgHZwK96qriUOCW2rPFmIuAEcVpdB7ZOUl4bV0uqTZOqCKjXEbzWyLx4RM8OcuS/
AXgRr/fuKR5zpTqZl7+QbtIrT3WdNskQW5ebykTotsg6vkc6ss9vVrDdTYNo4R2Z
rdkDKlbAYF/Q83+ZE9vIoHoZ6+Yv/ldAhh5SLrwQCki650rC5hN/CBIPwRGaBW57
pACIauhiNCItyPlZJLHXjdSxI0n+w8di0wanM2oZdZBX6/CFW+S0gv8LEsiskvgd
3QKsafnsXfSju1sKcP4PK9L5TqjN2H58CPZbK7g4wTz5frTAdNBjmFsgp7lZ75bd
AbWKKifqSlQHJqrnAYx1Nvf6d+SiGP6/J+r6J1bTrVHhH0tB0g++9kBScsZLTEV8
BeS4uyhKc8IdeMKQCw8V2SJ46KuzOG/PjjdoghUpJb0+qwA8p2ZTAFDKhH5UTkat
o1znCB5ebVZi2ojSFrF9epuStplaMJ+0C5tlLWpdD+95AFLJK6F7oTvdbo/ZKhfQ
HcRWP//4ncyAPWm5cArgm1e30hm6//R1VpadQk/03QmxBuyDSW+jJaVGPfRwKoIl
/SK54hBTMM0apywCbwxpqOenwgoI8UAcwLESxtSbZ28/lc/sVVUXXiuRo26L/PNE
6jpLXN7jSQMFI3AJVlhCDDdSc0J5rubQkzcLKVYUpF+lTtjJ/4rKC6Js3PR2pWI7
BGIS4ndfRjN6Y+WXbsLWEZO/viFPLmRV0ISD6ZxN+104YG+Ijsb3/g1Iey4/myCo
vFaHMDQ3g4jre12/ZOfBO15bRGRwL/GsIZyD537DVIL4flxjWYvqUsYw/HKSu5WE
IV9YGfiK0kyJU1Mp5iv4dmcGJmC4IdD1I/uUvEpUmDr8vZDgWYMD+lZzevmoQV3W
Z5ukJR47qeVXBIATn129xBRZcqQqLC0wFKI2UQ5G9LY/mDBDsrT+nZ2jbgcrAV9P
5ipDLJOCtIdEgeyQhdeiISb2a7I7h5j8UTqGHv0vqHsLYi0hB4GRoLMpZC1F1oH0
+YmzaIjb/PI5/0oR1QWbmDAWqaCAmiiMBJL7vMlWPyZLHTv+ch5dWTadJc+eFZwr
0knm26syDHblNNVDEAMH9c/dzmSGPeg80y1g02iOdCjIhR1K9zqyhLu5Nw6wFAl/
uefZwxApyQqZZTyPHs8Vl8CkBYuoNsqdN5sc1JyeEbKM208j5Kb8B0NpL4pZTyGO
AuB2AHNGfgeduHIYN63aT/RvUn+DM3xszE4F0qIF1B/VfK8unqIFT40PsAfvzrua
eY/ju1H+WfLfHMF8HDl8FDSaqizEaY1l/W1Nm7SF29i2UnJfbI49WNptgV0pdWiN
UVrtKs5alJ//4J9GEyA5njgSofAP+/FjVQvbjTaq8MSUl1eEE9AmpNbEIOszGOwU
iJiqm3TdpJC3MF782KJsPztpoI9GtLRgCoz004vkVTfEsiMS9GyHydwQw9gl7iRY
pUmNIN/ogBk1nBF+O/b1QB9Iv8CswWN50RFsXhspFCWJ+06cgE94hbC/2Pzc0OMA
ycQf0h7qm2fy0cYuKxvLxPJf3VnBoZt4VhuuXenMt6GLl9+RySPQ5V/wm4330Acz
Ak2Eynfky7R7DUwVZzxa31j+YMnJ7wj30iMNj25z7Ek8MNOTFamEKw40OIj7lLqL
jGaSH/f8MXxCEBqVHxwgNSRlHDQCGd5nz3KB9NBRSx9vUcnnfM53UTOnCTvGT/Mh
appVWJMNITZN3sEyvAOhWIssGtMEci6x57UL31z/lXi6YUrr8jBTLMEfm+JkaX09
FIaRx8HnxsjW3M0mEgK/U5PT35qV8/RCADw+OP2/y5Y9p/pnQ3Ib2ZWXxPL3BHZ7
XDyiMlDiObSts+VMMBwt+eeRFRH32o5U9VTJVAepLlWcnyQC1sY0ScTJo2C2kKB4
lJiBGdaOXV+CVyxfdAV8XeEHCtUNjbXkpuFPF6B0fIwa1kvLtMvwkG7j57mxbfrj
TBrslSWr+OwhbkhuJs4St2Xtd23ikMGkH6wnYILjMpyQ9E2xGEymHSfcz/6cVcen
tw/lR2UqMIrLsZOvM1o2DWwSE6q/R1r0tB/hO/n6mt4G/IZ+0ZFpyiTVMGE+3K2Z
x9xylmuAmLP8g9rr3t21CsKomRrP5slLqvX2rJHzKd2OD7l/6FRyD0VrzNHQx2uw
YO14SkyqIliZKpeGHm+q/hlwIOZ+SJ/mO9m9Oz2UYhFCrETwDZlQ9G2tHHm5M34Y
sWgphDQoN+yjH8prFzGIySoFTm/BS+EJ04ISERysg9jjVqXrZs4NkytE/VMgr0zV
1Jv9PEQgX9Ff8x1fkIcVajr56Iz8eF9vEp6OHSZsWRW7ZblIdZW+f07SZnND3NVb
xhnpJ/yuB9P843YF/vJnOVdx1jSpVuqFjpqy9yvNYl4s73W16Rzu7HMSdvga8rd8
LE8PkUh2hvBRMnNS42lxqdQlwNtU+e/aEG3YT7YF+DVSp/l5pXeK4qGWy6Ugq1TG
uIRcz62Lc8rsq9mSl3vVOl1F4D6O2ZlMnWEZbdP4cioaRwODXFHOAtVdsZ+1W5r9
NDXCy85mHABzXRg/JbGfQElYqRxpdc9CCyU5oqYvwJqCpnKlBM3TZ3Pwin3EFiZR
8k6hD5ti9iqz0okdSBkx3ugbLiY7OQPEgG7ilqEezNRj2Zf3TAcFTvhxTJKQYgZA
meQrJLMQ5HPN2gJvIG91yFBUafK2K2ICw+MeimwjO1pQeG+VxiGMUw5Ah0EtMKJW
zdwak1fYA+4arTF8OxmUJzFqZVjL+9sASsA7ys/7IH346JfDgP/4lGlrgrbT1qHi
BweFwoW7xCegn0BeGDevu1AC6g2ARfCbmyMSqMcTSAc18HLlsuM8ItYZP24b79An
Bloiz7TT/6Wduuy9Icfq3ikbB6TkMme4SVDrw8FNmtz/sBGYv41gb89sCuFxnWLY
OgWUUvfS0VyIkbGaxNddHTpzF32NCKxynSkW+I97GNUOVKk0+TsSkCL6SVgr4zi7
4X768fxuH8ZmCwbTwhuM5YxiyVygURv5GeIn69OXJPn+n5B+auENat1w+9u1DvvI
yU34waRD5+iFOzo0pzR/9PoYph8aLKw3barMMeZl8wg7dmCZZdhKxBThwQKkQ2sv
FJijX3yAUZdNmIUGeI5tIoUar4XFHBS0rF2CQy7r8usQfea4jDf2p8vRG6kSp4FC
/OUBRGR9cdfsO/AV8O8l09x0WkUT1bT82QpX66/f2uCAtuZnTJxtKsiXCYjT961D
7dSF5Za2ALNdvWGcM45d+SB98SmxBpAVgYfMi5F8LsneMN/rW3aKsBFg9Bg9kqc/
M7M12WRz76HpnfujS8+FZFnhovPlVBtXAtAeks0pbvDLcEtfYTPsILNJuVWYbchX
ONtXJvRY8WZzJ4ek/1HHbN2G4IGPRvJIMlxx3ji70cy0V6VyqCdMcLX665ccqCCk
xJo3aA/VBFxFlToqDiy38LOIOtotDcGsgZfQmGjvGnhlT3HwL9/dj1hcrLriM7NI
Bg8rcLDZvh6RWVBEO4QEbWHrQtvzJgLGCY/79jGixsvayw6AFO9c0jf/6A9WOrg4
aZtEdGTkgZrwPUx3A6wKKV5OcKT9M4HzMB+M8dtEY9Hhv/7JmXSCJOiTILu5N+q4
1zj2c/lRH4NNWmmh5JMj6pYc9ihAq1IHJtmwWxBQmam/ZnT1kJmgBPltSLUPduTt
Fez0RH3a9vzvLQGDAYlV4XohWlLoRZynPHWDFE381gfE+vdRi03E5RBEXHXYhW6c
0C9IRZjnhzUAc7ewGk/4m89xBEt6j39ORXzqJcO0ulJlg33VLjmfBBjZ12DOXlo/
y9yzQrYXtVD2UtrxrfzSLVEh3oaVc3Ck1pQoHhM9qJ9kdeFFHydcBSRi5qP2mEIs
bhQJY+XD2v28JIqMFkbKAefKwSa0turt/P4B4BHSbH7EXY9GAN8OfqpTG0K0CiXx
3XAsE02tv920QtcgX2pz019Vq9r0acN8AuFTa1xpht9RLT446zEdmQflojBiDhbw
vgaAtjjDxFo2ZYbwAAjwUpRsBYixX3u4/F2OhDQICWYW5G8oUtWj9Qzpljmey9q1
6kTGYysHMoGtrsr82h4hqZyyKWnOip3jtAfD5MoerzLnBUSNurFc4Y5cDpfGNTXN
S/x9ybDmzVpnqDIPlOiQ/gm2bkIdAquQ02/6cG7KM8oxwg9QpubuXBdfvVjSoOpU
gUY1QsxgIFjdz7KB0iVp7egOpLJB91n0MIDnSt8ITBEWgVzj4QMZVpYW2fvlWfIl
R9iagC7PBkq/Fd5do3QQiPcPLryfZhrdG4YBCOFhqp3sBnuVKVGJtEp3+5I+IiRT
/PEoi16camInVLw/s0GQsD1cjMmzucdo+/a+fXJGAEJHY007i0iC2YEO/ijMZTYj
L31eSAqrggPT4hQESgALcoRiu/EPnU2UJ5K4TnSaW2/3l36Mp8DYF4ew8364S1xk
Ljg2ze5ACkpjXP/Wui/c8heuMVn86K8YLCEFx9rG0Cxr/ytDtgZAHNY/cFgOlPEX
HeO7vHbU005mfafhaG/snlK/uOiqTpDt81HaSzlVEpqMOj8DZ0fwIl13OFysLePB
KCtyKI7PhBV4ktVULcaaV+tp9uVVRPYD6bjBmseqB/SH25th7IlCKdnF1xcSKPb7
rNxVVnYoRaAJ7NC0XIt88pqsmFepAdCjqEex0BB4TegNVQ79FFhOQHM6m47wnQI/
CzpW7iISAKx/btVZ9ylKDVUM3q5dYYE4rAojASW7gdDlC+qEz2Ezr/v8qL2oJ3cL
1XehDUNBYOBf7+ZtpbnJtxuAPrd2L/N/cwJ4GxaRWApXcxHop874EKtO4tgaqaeS
zxd2midrho05wnL3THvvyuuiJdfSKjy80anTddlT+WtSnc9rBktIzD5NtljcXZf0
yJQ/eHVTTB2FDzKeYnZmN3JhYu7uwdaYs0WsfbNo/RvqExxXPelPK6KJQIIYkf/h
1RIB8THEGB7rowaCodyhk9Lpdq7o55rcqU3EVwQ6a1rWk4dEGnFRirbHKXCICWpB
0ei7WMFGdrPHQDfoNy2YExgX52hTdNtt1jzTr4WYP7HChG+Aah9MZST7ayp8JXhg
Pxp9xK+Vnhxj6slK9lsQf0crOkGDGcx5la+QFAA8hc4TReiiCTZUxlzVMFBf0GvJ
zp0APTMO+j3LCwPAgNf5R8/MnC4yQG4OSoFf3hc6P5J6baHK6/vvRLVDFRuF4LwM
8V+F6BZ6HIOS4OpiICZNeO7peoI10d3sBABC+l76pcptsb7hZyj7buZdYccibStX
C/wfWHklouzJ63RC5p2ZSm6iiIJpJY05voRFEynviDJgxmVgHCYPaRzMjh1ixngI
BZgIaAy5yRLkUGJjUYrmgwN9aEB671oiciBXlgoKdrVAAN+reQnrM62C9lj/dqMt
1Oh6aufvpra5pPCAP4MFBKUxEcW+7uqEMJB9BpwBz4O0wutYt5vBfIlVDQFxaCOn
FAp3En9aa2HMqV/p1lgzo66oTLn6KgJbAymXHyTKmcTGcbgtUDB3amuwErPHF5CZ
tIbBW85xa0ReYeGNbx3XV1cOJdpr4mBpRTZR9TI0O9mnAoPRbC4EtC7g/2Px+woY
xRaNjdPfh5LBkmxJdsMZN2hx5F8tlK+GZdRKNgA+Hu7kCe6eMPF09EHYSFIgeJ0w
/07WUg20t+z6eM2nbCRpxiF0eZS3HIDw7+hTwm0exRcXSzUGOfbHsIE1hRNysTji
WcmeoBxdz3lUEDclIPOh4T2qELhlbX9YylASxKPZbJ4jLoC4BVUluTcIkG2F4CAB
sQY7X6SVz3VDe36I4n2QLxVkze+iB43hV9PyRO1ZVzOpCtIhse2690xjnZBnyGSi
PxcQMAgDT+mnB82bbLpHm4vtlMnfg+j6P4/hEZHVugr1gzEiqhLjxTUfR72UECfW
tNozUuEceOrfz9BEsqLMQQjXnBEEL4ApU7EWHXX4Xn/cbbeBFDkjS8FDc7SEhRwc
Wzgg0DfKVSq72OxOUW4XC1O4L9pxjF5C1lzLwZICdTd/EnUZnMZHnLvsSnZnu3rx
4KROfe7hSTBRMZJItnM1vdid85DYjcMLIj6XAwMvO9Y+6mbmGVWgqyfoqx7YCUE8
nlJSjRE8WXdbGzMQMah/Lnh7MYiqvkUVniQVGVZmjh4w2mPAmocxjeP/PcXRr4H0
hXKduCB7sBa9bOQFV8kVyxzsKm6aAYoCCfBrhhiTNJmu4y08yADMZNhzCrkGISpr
GfKtAaQ2y+d7Q2fpXPNl7qc2pdTLrIOJnQ34x4ijojPFyMJvYOf9ZgWTFsE2Gz+y
2ElujsSMiR3wBroCV9QIodc+3hg8c4Eh/KxqzAl2yBkw7FW414TVQTCsOgOzNc8U
J7ClE3I99B10bIbA8kETPRhCr2fI+N6sNojGWsK/52yzzKRq6BarC2q/1PPUQABx
C65pphm/tjqOAJjG8PGa3W+Ma6xBuwaKzeJoExl+EVixzU+W3946aKRZ3XTVrqhH
aUIhzTfGggWEgAJ8NzRpWjylpdefytO8c4u3RCUA2a4eWj7Al5b7U/p7lmtTnNpv
ogejYiL8+7vIP5C9WlTMVvUB4FHl/gJmbx9JFsdfoP9wkWHT+vCiSuKsFJ5QTPI8
Vf3Lem53wwStsVdAfpvGuBdhneaGoLgRRHCI+LlDdR/uEPvp0p0tferz3y/5NB1P
Cl6nTjNewOaDh0RCTL4hqWw1C5lp9S41u7WrLYax2Ho8jByBqY+BPwLs2QFyFyG5
uPYjmKotFpPTAynaufc3OIGow6AA7fSzTvQFXg8MZJzvKNwXJJXMHb7tUEPRjWyg
LphPkKDJH3iQ8StGEDRLmYxvJ/Ik5mvZAmmLGi2vuF/WT6AMd59DOLzS9ojemanj
vezCo7IE6v+whv1IeYWTdVtOVF1998tTrpCTLepXiKCob+cxx63vRskswCorgcEg
5Zmjd6Wq5FJLaOKAggsGc5d7cWss1OUEZbLQZcDxwJ27bZZdYxnZVgo6XqbW7AZk
u6m4D2zmNiuQk49QCHcFjyl8dmjAMDVbb7BYSTIRHERhR6mIbqw6YJE60/i779qf
loa0BvdR0Lryn5vJlEFmj/dUaGF1twZ0WGp98HrgvhxZcCgh+bn6drmRvplfT6bd
TDFwW06O3c2bN9+BjZ0qlHJBkmks36v6pB8OrcqqJwsbthYQJ8VsKL7jggq1bhSf
XuYOZZDDKWBoRwSkqbLXo94XqMx7+RMz1oERu2aseJoAwyBV1a9vLYTAz5Ac2s5B
vpegTh+lR88WgZRSZSuxx1iham0jtqrpNtiXIukFSwxgrROyY4EBTGv2tGJnmpcL
0JeGc8VxajCxHRNvWxNCP5yFhHb+31RX4lAWOqcvApwrx+24MrMTWWCGdzhwmWRX
2rCzCAtYPbWmpIJAZZHJxz1JNuQho1YQzZU+h4nlLZyKEVlXh9P7NoyQPE8N/Jnr
GfoLrIiLTJmWRdTQU7NbbZdVsDtCB5EwAVb7b7w2MVP39xvDhJ7u1RRsHgcJevXx
7K05Yk8S424Za0QpVAadHhZSsI+T7lxVqsCMgCNFTxc1E2EjQU0IeG90n9mnuxJW
g+gBG0+C1y0jBeiK2WWUa8Ewd01Uz3P45YrTt8GJupYAPhz1m7FNGCvU5/Fg7mah
Dg6/pVgblYk5BqTuTtl15AKs+0Mhc4P0GyO5JHKp6DbC66pFaKuoTWKxD1N2V4q9
Peiexod7HPa/wkwLERBzOk8s1Rzx10s1FTqr4HBjT3+EkOG+faRq2RFvwiSyHmOK
g6dGIjXgs/5u7EDow1cmkjsOcquFdkIKeFgEwOd1wsqXCt7lzmZInrra4+rSgOsb
Jy+Ml2vt1qu0+umrAk8FgJEQog55jzm1f9JA9ySEtru8jbR41vtbS7NoxHeXnUyX
jyBGACcz/ep5O38KrtAuDSMWZwZm0kdkROfqQbDh1F9Vp+BbR6iFmNPTNPHWJxhR
hD5Es41RbCpI1dvNyZJErV29DsZWDpbchCGaVK01t1+fjxTtOAdwbVEnCA98bg9l
uV/sDiORJXCHel325Dcv3rQ4AoibeMgknT5+YyGh97j0sF33kQ7qFuAw2/aD2lTL
OdohHhwsidR40ujQ+uuadtmg8CSaVILMYPJWFSNs6NVmIBkZGsr/xZ/G3egjpCKz
KdcWCLbYgRgyBrpVgJno47vhVpM9FPv3pzdD+WOM+MbB+R3gWUbefsAwKAZe1JxD
iRGJrYi5mGk/kmFGGk6hwzUNfdt5ltSdN3MnHx5/549D6FybSeFhIKJ7fAkt6poA
UZFVm728U9Jnmnpbq287R74p8uZHy6b6Lv3qXAH5qH7K0JzL7hlMPsclcmEjcltm
S6AhorxFDzcpEIxtJvjEOzIZgF5Zv9bPKBTjU/siIDOLReUyPwDYZIuoLi9Gm201
COK1U0xZwi117IRtgg9Jlc/E3lojT9vhA/tN2+GA4Tl8bwfppMIwLgc5bLPi8TID
aSw0ZZFE/RMtmcy9EAYuAsTQfiqbxR+b7QIfBvEaUUD/MlGGkl0Bh+mhP8N4z+6I
Jj3hdRGUpgbjaYhieZsU6iPEqefgkt3r0RQsb9zFWlis2JxGTqqD1drtkq1xcvf7
UxrUOBZURdm28HDOusvb+hf+3dMvz3AvOJkfelVtC/q4aBYHkFCBWNpXWYk3GmsG
tM1uzBTfkqcV7kVk084npCZ/hh5zP2CXPxWYpaVkftuBFiFNg4frMawiVDgB9JF1
cYtPrVD6jebhzxXac0CEBH/Ix4z7snV1o0zWN7YKYw9OpF0AYYtcuwJs5bCF9DLn
r0NzUENCsz/6f7ARGDSEGI9Fy57YR3IgXnMKKYQmTt3Pfhcmmcefci59klnjB+NI
BrQEcM8wH/mpomoFo/jGYxnIJrdIFbLAwiIDw0a+NADSkHFUmC+x4jm93ZOrcyL8
K5fLnYcnt1II+9jFQachCrMsgPtjFQ4eHYAfh22YMX336UNGcZJIqaUhsbKR4rAY
LymfOB/UzYwLhavH0tbl1dtprbNse79Wq7gyGgH/nxmvCGfpuXSWNAPTeqkaCz0S
3q2qzLvINMjA/gZcc6FFBEbKgYI+HZuQp6XHR0sl/LPg/7T/qeLppeNfopu+rE00
Sk26QuatEwNgegzqQUiGMJ8YRo/IpngxnsWZ4QYCh4BtulB5MZgH971GaS83XJDF
sPhPZkaUXXsqTWTSzPUgZ+acb3j7aThyhMXEvosVi5lRr9JlmgOKku/FRH4v4HoO
pRuM6D4NY1MWMXAw71jSlxGuYCbwKlQosbqD41HvLNUfFC9YBWNE439m3P3JmVNS
jC6LG8C7SFDx31s6gfzEIwuewVRRtgxMvw5Hi+No2dDMMCjohfbOqnO7FXm6mYiX
7YKmD05wtcfaglTlsXzTvNdQur0vbWr1SL5iMxRjT+QbrYnyEdpUlpm1mJLQ9m6s
EzyfB1pAabyk4nnx1xlYyY8An3NeatSYxC4X33ROfZEfhG5ogQOrXIHKKpP17ANw
BO2W+miOwDT/nORDJjk7aA5rda5ogoDvV6rnLOtdBZFOp24qL2T+Q0ubGEZkLD4D
qD9/KEdBm6ce428uIGqgm0BTFeN99krnoJXC0hVID+bODSzcoO+8vrtmRg+0lthw
HAqzpYnzlgOOY/6bT4vpXIzIRuNuTOTDdhujiHwicfMpWgDa6D+S1+AMSYMQ+BcC
pUzic68RjSSugDXuKvsKYVVO3PcmyeZIOrNp8ZBsM6Extj19TyaYMAZny6SllUFz
nMBgnTSy8OTVOIehWOdzyfm9myvFKfyv660g7Kd3FoGIE+rQBDACZdYrHZJwbnIo
7eROsuNFiQR/8LSUf6QAD1X841DBccXJl96qYMZ9XXk4638h470m4jsrmFD7tGYB
/GL3fLyu4JX/Otqobogwl1RDBq2HqHEx374iQxUDEIDD0WAT0KjBV27OGmFgWBLp
g8/tNTE4fPXiBDdYbbDemi0IRSAYv3/xgbanC3lnIWhaCHgqCHIzA4OvKLprL9zH
it7l7s5vA6+/DatvQdakUAaxg4pfpeKcgyj5pIT3saMzrRYMkiesd757pQKSVEcE
H9EnjZX/XGAqSp/59TBHoqf0ObL4vtQaH3sXG02N/SQ1mD2h0SHyt4BTnTWKg5Cg
41TcgdWSg7MyohJsVqIJAKYzTqxI+LArp9dlosInOynt4DyuE5k03L8TJnaQJv/F
U7bMJ/u/l2a6w5LPR+dGk5zB/JdmFW6dld/uWvSOO8HEVLj0dGFfnr2lqDNepUGG
jJ0tHk8yDfUNhWTuMd1wRHgHQnO68aoRwRps098D1bNS+dwfHDO6hiT+GL4pUs6D
djRBY+p2I8q2Pj9PIegxVWDnmCcXelM79QUa8oYlgwiyie6aQBlAQp10yxZvNuhn
tm90gcwsXZYTx6RQNfoJA7TkqsSEEh070E1fx/9IaH2qDpcOdxv8qxdsqRMUNDdX
JTxL0pQvhE/DU2x8NEhG8Tn5XXwX3D6rQ5ZwIyVmQCy3oEpAGWdXDmxS8ENOT25y
lMnsof7GYQHW9hJpbBt4BHOfpiB6BCZ3YD0Bdnz5Cg+IkUYltuCIRmstaKuJ4Vk3
8mWwZbpFUOln+UXDgk4dtaeqSXK7zw7uls4ls7FbgvxN46C6/XXzR1s27ppnhNpl
JHdXQ/sv14dVnHSIHL1gyie75ksm9dUzYg9rt1McxJvuTmBDSDXSQtbwaa/DUfXz
MN9aCJuJQM26C/gG9QQh1RCWuiu4PlXKhr1ROD9SEuoGgnGVXics6mFC60ynRO3K
wXFb4HCCvtLzktgFxu1JqRnlloVPh0FABZINtPclS1VDUFP/reM9mJU2iKOiuA9g
pE6gYD4yDUgF+7aZrBQNfaZ+utXlUxmoYFJ6cKwCrdarQ18aE7bdRyQhjHtDgLsv
mx2ejWEkVlMiYjH03Yuf8n2D+brNjjtEPzBQVbxVeImmuAtdqUAibcKwYxIaTfJl
VRSzBby8jVZfKuKSyAoE78zTQE+yUFr6zrYiysbFR6aLFQpM/JPJWhTmoHJ+qh3m
xXTha2W0hg/au+3Vd8KfRkqoJ1CLHOo7znb+jgvYXYkynfw8gPHgR2ncLTpJPVXu
8UKWLU/Qg3P9rJvVxqV+89fMKELejT498IwD2HJ/sWHCgZKA+OVxXDQX/QGD4d5w
4AU10K8m8o4bs52l7rjw4ubMGAVC6hP7oEQFy7Kfuf9Ec7unDPmBJeRBOfA9J+VY
HNofHNNhe/7XyOgskybssrNz6W3Qd0QYio3ao5y0OtMIqmt197eRWXYre1HuoxP2
IOgNGZ32Sfu1SErXBW2z42sdt6nAARVx4o0Mt61yew6swwwAKMUE+MqEGH+g41u+
NHKld7hJr6oVBwth4x8CJSQBUGP9e2aDRYksUPhjjnvN8fYQ9IkOyCa7UTJDpzqP
Wh7TRIcSlU4oxzd68/J+Re/gkcF3q3CqlIYldX47XSQAv/UUpuwy6Y0CWPx/XLZH
p3IQDwEn+pV9qCIFvr8Ni5r4DubQDbnUrivkQzKfLgHP0+sB8QLXofhAFvzEFDAr
IudNc03pf2lvsetLKIqND204obAvARA7QPDpsuwgc5TY8xdARUD8GGlQNQCIIbQZ
BCGm570/vecLvuXqTSMWprnU39hO1SqrjMgUGoMFmXbeJMfZkCmJccHPGAKvoZi4
BtBHp7URyU4MoCLBTEZQ5WsN2Ea+4ovpDKayGXNlqyNdxDf2Dqu1ydcQlf56PqdP
uOp1dRhb7zi41MDsW0AWBPPbSHgbFhY8g/dShfm+Gb3NpfV10rS+A9RRLb9Ww8cO
5POLfGJLxFUr3plSpgTQUwWg/pHi17AcDdqpNHWUPJ1H+QfCG9PCstcCS5A1Q5hf
Edps6T3a/4B00/2kILdz9npgARWRUL/HMIymMqqbM1BeFxNe3zvqkVBSBfMDdTJ7
u5HdoBgNH9bDZo0mUztz/PNmMCbCWbTg+TXnH/mVMTx73WMdv1uy6jnyvhBxzrwy
ji+0QSQaSkRB7IIfp4sFQZrswCe+l3Pn9AsKmCphKXCpaqJsOuU6yP602mxg1aCn
q+9MwgNmmilnxRQafxuAd/vd3Qx7RjdzovMz7PrIlPe3XzEtTQDsBfcgWg4IvQAq
lpQB56shyK/cknWoL7G8tlYFAtNIBqE/R3PDcbXoL8GRdAGX1VEP0ZkcydkWb03W
2n2rdOqLagCRCYxxCbrlKbrTTEfLxvs24F8apcJILs2kiQvmxbqCGS9Mt11lZtS2
Z4/I2Wljya/vFtTtTgjWBTK5JXbynqkhbfUqm2cUTSxwBrfzmInJikUvUJ23qWF+
cAUbfL8Ati3SkZAALPix96HNWD3LJWXinaapiwTwLIK6L46qWJuI22LiRdtjx9tx
JGqOxudUfM9Zxrnwfd7bURP3HJe65jJuq1T5aZf2V9efcX1ptJbKe1QLHyqC8QT6
aifBapvFFsWrlxsB/fokLGjMZcLPraUJBJDf4+UYnxCwOgmk0Q/HGAEfYAlocfxV
lsCsFnsEms3+VQtRHXL6QfGwTPUBaIAu4DeG6G2AML5ycqSwCgP3M5bIjWyu/5ON
VRBXoMhUltc0o5TaEa3pR/cdkmuK1cCUSWZ7KZWK+rlHBWaq+NXHJ4HNRJycP2M2
91ZwyOwCbsrVAu2XHncZMvNYzRjxGx2Rkpq6wgX5SPP9xkxmWDF5KGOiZmywBXO6
InEY5NH37rlxDFnvGaSEDkwkZwlgBY2bST8jzrWOLZDVynlhoeek/7w3qe65Fklf
sIgQV/sldrvvgR8/lhI0DPLzn/HyNBhJ8M1MkLsSdPRHGliMafl197Pm+/OpqSgY
XKCo9JWvnH0RkJjRmYCjSXzD5lIR5Eo5/+hg3AF77Hu43IdLw8KxrIww0qnYvIq5
WAttmNEWPqBR7cnioKgyzeUOwDhI+4YCM8DMTLUvmx0/A2VnuBRzwPxDyuHIq4Po
pMvKYJodyPsctoEhgtGyFT1JpDNuQO50yoIRg9VeV+7UWpUdyjFachKK3lPx91Zq
4GtEJ0YiEwwtSOM888uftAR81JfHGJVAr+n2DPa14xyOdZVhRhrxaSzrpeO+6OBQ
yBUgoiYrtJQoYFVafo0wPRdAuPhPjmM6YOqgLsazVEjdrwR+Hu53RpZBQ3qO+wa4
Gn57kIfg/gyKH6SRstHNjifaMfB45GvB3jvvl7L/Ip2IOpTwRGysEJh9ybT0QS7Q
Z5S51wA4wxygVZE6AHfVlFn1aWGbYhyDE+90xSgvU4CEuonLQxtSdCfWt7OWSG+m
OFLqGbjP3ntfEXQ8BnQBdGkkmkQCYmy0QzHK0rADahAV4SJugm3mSpsbt6UKIIIl
9f7CEN0er2EMk1eRGa8QsdSMgXXS//+xQbz27tl97LW0bh1+SuexdVG6uOlVuNEE
a7tFYyPXL7ZV7YxAsGVoH0dg9eJ33nous1G5jGfjW26VH4W4FRWJGEsvkMXSwTjq
G7SQlz2aSsXdO3X0JrLO112pVRHLX96vo8/h0I8t65ezh6CA1oYZbOUN3ofxCkCr
lgKEJbxEFLwswH+nCbYBZslqaq856jLfkDgpXd29puENU3yogTsaNz7BPRW5C6Mo
M1G45CbRIaSlUJMDLmCVZjzlZ+rbCGz3BR2YhEoDi9FhAWyLpsWjRYLkHOdf8I9D
DWG8AfEfwkBNL767EWxRYynxUcAUOHTe4BInAdgFD+HpHRR6tQc3Q6g3bNzPR/o2
6pehpBFbSFTSvzNT18Fp/wEAO5dNSEpEi6IbauHttxTI10Ur5hMsyASNq96k3dr/
IlunNSmykhKqVsfQFxqm6fHPqtZzPhjQpH5wK5HXfzh1P1/FCKzmwCceNti7k9XB
NygTOwwEInic/x7KsqCEL6yvqwYFmhW/qUhxpU9m0CgwauVI2f+r3cnSZihp06gW
Frth5F1wWuXoRUXXhtzpCeUlpEr24gbzUsLuFQ5mSr5MfZqjM7w/najgfSMHONhO
p0CJmUOTz/atLrogcg9AzgcNiV3nu0Xukr0VE72VQ8t1i4eg7Sh0oy/Z/LZRO7V0
WuDg5RV6TFLYA5csUcPPbsKdI+jcBMgM1erhBh2wULXbZ3joYVBAPWfkqr6uwgD4
M/PHXpFro7Ku5oaRFjSx/mF61zU9kWftTCItMDslGzyxmbcO8BQ5aHvSVsFWv6Wj
EWzIeSLnmOR6J5BxOTSgZcbtZ8eq7G2VvWJgmL0nvz+nLabguVQLtNN7Wu2DxL2E
eIoa7DRp62VpBbB/x9HhbaNCIiUbX4aAdw7q0OOg0U+yj+qMly5LErYoXoXUVa3I
1ZRPepFzX/ZGEiiJCMuOdtMHxq2Jb7z/Bw7ZFhkxQ74SlE8DOeOzHZUCExK2GRNB
se1gAsAzw5Xs0i+XxCuUEy/Mjbs1ncnzF82H/nU0N8SITjqKYMw4qUFeJVjQG/zy
ho2SppSu2Sy2tXNRZAj308H+FZucwE8OFEQQgkjnoliLIW9Va0NV0p9udtdCuhlv
txD/uEXieyV/lQShX1Phvfbr9UwYrn1Fw3VDgdf06hu0syCxVsZu8oizH9Uh2nVn
XJpVJqMSiHv5P1d1oBtOqGkKYb37J7TDwtfahJ0IB3cLG4gSQaSBd2VELVACC6TE
wJqhxiTLBA3Kaby5S3uVJIPw6u5gSuZpUH1S6L1uFBUyjtGafvqzsvN6ZeCgSbfT
eKY+K0/cvMJMkLaG8XEWi72sMFli68F8N1d2moL/NKG+cskKFR0mtW0ThvctolVB
/diGdiSYx8A8QdCLTb1tJdFsOFOBNxtg74SEw4saPyBRjFCSK7cSDdCrmQ7ltH8u
+g1q2wAyKxqVqG3mm2Dh+Qf9zMobT1O5UCJ0giM/Nm5nuyKk8l3JJP/9UcH/S9Sk
oudoYlKHhCdVoVfScVRjZYvZN0oZ1wECxu6rw9zJqWdFrskSyxHRXCdlMvIXdD8f
0j3OFCY49p+W5cHOuPZUnpapZ1Cv8fkbjNNqGG48TxQI6z+YC5YUG2kPP8CHlpOj
T+JNLkUUfCJKNc7yRF+ZHyvSKHTZmkSca0HH0S7jxcBBRhVtzy6KfjRWEN9yo2I8
phYYtFaoOhtO21kxpBNEaXLpyuaZFlbb5kaVjDVxTjdurMMqigFw05gLs2DcALu2
o7H9QU+5y80uw2n7v7LE9/sTpypfbdNl646QbEAvb+nXHzRLVXQIE/UjyDnZFSxc
ovJTQFfUzUH3zxNuiuUW9o4SeQ96umQ+N7wPWyWx5+YCRpKW9bypP+vtx9/4LqS1
Mq6LgrzY2RnxfI8O9juBp4uzUoGSwtEonYpmnl2eb+P279MD8lCeegIdxMDEMZE3
0KXSg8CaHrIRvmwPKGukLImBvuga871DZCXnON9viMO/8ZS+WCYucUQxsDXhSvwr
Me4fTSAnQnJaxK3JKOf5KmHxuhOuErO04x6xNEtYqkKoTjDk/lwJulxBTrQQobjd
6bKY3YMFzSb59MbKGFaVt80YX49KHxVL/WCvg95k/bnNC8RlwTHFUgIacjQrGEvM
3DACFBNdfcC8dbKXj3sR9K7x0386r7wbvPXUrRMt4jTp9+sNPHyHL0H9T6z4tFgm
Hb8ebDHt5OJ9Syb4zDmY2+IwEi+rFzsWHiOGwDz3/H2+GWr1OXphlnvYEf2pDKh8
PmMKDO/exilKqx9W05eGvsUXohF+2PWOnfNxmxP07nZu/9K7Gk1EU8llMGYI+nnA
P0lwwNBaasaOB7/ZpR/2VQ6gxoBERwoIRZEYtmJ4a+COKHues2zGue8Ji1t9AGqd
X4FTL4dpdhbXFt+IIBmi0XDAiV9LCPEXESPzGZ3kc2BR36iU6VozI36FIrqF4GAT
wa4is0ts/ZrJSlVnGfPyk5jey+2Vu1/wA0/gfDjxa4HybJqd9L7l+tMiaBwkWR2+
g4yRJd6z2hA43+DYIUAZZYRfteAElorTWIn0WTAyE7KYIIso7dTp8tVqlHkpeGMH
BApYXLxn9J1ZpI+v5yQY/rRLiYBAAyAHSrvMdDPmg383h79F0dJvy0ajyx9ZA5gT
Y66TRd6tdEfxYITup138TinrGL7dfO5Ep68VpDLrlRa+GcNYQoLpiXB0E3A6owvR
Th9L+sWtZElfPHICZWil6dHan0LoTDiJ1D3G97bj4asGe0E6NC9DESaDT4WQIanK
vmNbZ8ZU3jS+9IDG71jMcqy/Fp1uNB/2/yBZ0nPJTpDiYir2sbHRGLoTqS9UoGOQ
UkUa6rNY8rfYxFuQsz7uFGMbW4UBXU/XHg992LXH/Wfr6yDrzCXdrHtxE8tSDczH
CGZrnBbQFJK8DP+dHZAE+vq7Ag4lN4vC+mSiD9bmkZfRHKoPLFN3ehCIugcM1gOC
r5B5TJQr+O7GtQyIhgkaT36FB+fF+hAiPiKYsyEml0GXWYZq7D+FrWiE28+68a8w
zBNK4MIyO0X9KkwTRVLpf9Gp5Bb64ZflykJX5IMZ/x0rf6/BV4xcWSGQvIiF8Wqw
jY7nOWcCZd5SDgQMuHtQX0xZYuba1l8aw45iUTN2kwp01pVbqKY4pUMpvaAFeRD6
pwVpnEPuoFFvbpUNkuM1raUU1SuScbWAlaCZFzovlrhqlfcsON3mG2+W8oRsSFLe
lLqLpP5fAUvCtFra+MwKyWg2q72xrize5j4r8FhyN6HNxLXrPmOUwweZSEnqW2VG
EMb2LcpTXTXAPIldNRK/WgUCahkH5ZesyMQEUiO63cjRii7fFN3AEHKED93jwoGO
6BCySJRqsSxzX6GJv8tIUhaYR14juuq/+ZqRxN9ih1SERwbp+lnRwiget1XifRCR
u0Ye+TFLE3zLJh90SbN+vlsgXwtbwcTSbUyeFNnzd4D2hqHI8plF0T26xXVTYnRC
DQqIstqq2HhJ7FXIhbJTGNScew9+Zlc5JwG7zR3Yb3w4yu4+PRMk/rzZpjAbAeF0
qoABWqFYHAJ1kIO6aPjX66E3t4/PHM9gCwIDbrVlGTtliVTf0V6xNmd7uWu1bzh3
EJrI+Xqe58AjO/VBI4GR6skPmMsJHbU0HT5PVW+nnRCx+jkDKR3MtZPJxD5XA8Hq
FhCVkIHmQs7oYMER968J+6AZHclqOD7HD6V95445oa1qOimFDLz80gpi9BXRj4+8
D7J+ST1dnB5NtLEGy1N9DWevMUuXvRdtXESY8FMmfeEN6U3MbqpVesKlWJMqn98r
aBEcEHouKGImTsQFI0xq2KRQc5U3xeOX/pe8BRS8T09Vg1Q6WBqF+DDP9D2uSXAz
67vnyNb5ixwPiRxKNZjn2uf4kKy1Of8TZI2wcrP8ZVauhJwFRp4nQT4OaWxiq3PV
PxuJW1J2X19NQLRtJKppD1dAd8PASVyQACfcQlhdAH9eGBodeaq4hLBqK0ZmdS7g
ESCQgM8Tl5zb3VQ303NdGLxNWnjb+bnfstTykzJAL/GVXliq0S9Di7vpmhVWUeFC
WEhnGj2Y4MekOSiy75G9q7Hcljw12xXLMZpF2pr9A96ohV+ide2BBt8vU075oL3D
fgEizAjjKWFHlPPTpBF8E30wN3g04CqHlTMy2dlWK0pWexYPjT0U53h8VrDHzI47
EP/F2mqf9WI2fkdaBuRm6HrDq4hVSyRw3819HasYYv2uhiDdZE2+P+ZNAF2GHJYB
8+Incnbp1ngPJNUkc9XQmvwvFZcSoVAsQLpt4T2MZlFFVJpjzFY4SxrLjyDeY+7S
MjINg+EnSAgrosyLp6gfQnMEM/0bT/qOK8z5Randfn+E34vJTvXCL5Kbz+jguT3g
B/NzTes0b9VNJ0M3XHYxgPERDyWE9Hi7+oicxP5d+IHwehEPZaBrntZ0YIJtDxzq
GMltA3jPINyAgmQT5u0zBJaLa3knwspnPeTDUpJl+qdB8lLNE6hpgybmqOOLUnFF
4bDwFmMaci8I0I5UkUl2UMZ/qU9g1szP3bk3wrTKTvmaDePTJb2ehJqnPkVmCRjZ
ZlwG4f99fRTn7AcVQd9xuofJaxoL1VR0EmQAJTCaCebz9kYllDFhCjkJtZOxBqdL
EXFEgc2yLIE31ZyNufdS9Nr7VGlpxkaSCkT51SaK9O6Zj9Xm3apVlz9VRX0XGCaO
8yQVZuI2t3Z1kyN7ozRyChmbeTxeooywzCGfTbSuXr2rApPLIs256f9BhB8H64lP
0aqfz/sRBsijeO6nhNEVb9VWpZW8xOAFVGxoQCT8jvWAPfP0b3nczA9kSdGszxiP
tgy9O53lZctdBZreyWQnc+GtWQtudXC2h0p0o9In0pEkGqYy/vdb82SnyP8bEPTi
GpIxlJhB7plbdwhJ+okJY0ZwQFhYffHixMotBEY2lcdBQ/tjSJ+BbNj2OdAARR+C
BjNpxZMTrYA3ViPiUrhXN9FmPFSo3SzSykFAaY6+fS7b3lBzyheC6vT7ElooYPVQ
yIdySOsG2X2KIwDXBNjn9flN9taF3DlJoHsp/vGxJaFPL06HJKbKA9g1qpq1Sd7l
pa2FIqLkdYBc1rYW9y20h+y6h9CZZQ5QAKMjqN83Z0ekQIlkHxzsuScaVpXG00IO
iao5kQzEJW1JAiigf33JizW8UZcrDmdPOsuk7YcYhmtyy7rzt3LKlB9XfrT9tEr3
okQKJgjgiQSYpaD/KeuInYfrwsez9O1WdUmBzGHTwEH0ctDxQ7MbrxAupaP66ZGI
g7GhQuIlANrgfBGd5sQspeYDviI+A/wUnfzPhZsg7b3Fc+U1g0x/Wli4hs4BUGMM
GQVGWsJCv3j/biKItpMw4TmyO2o/5iBzSBAF7Lsfd2zTY2T6obDrh6FFQqURSpHS
HnsxYiw7KbOwdtGk6Bf+g05uTu34myLGj2F/LALRvtVNfo7vfIY+OYqPtnbgiSgg
SMTqYR/97x8JdoXPMX/RDvb7j03BIMNLvshdEwiU5Nq2XvLL7AfzLUPzI38XvvBS
p/2YPbggjPdYk6wixxRL/tmFYaxTavdP0iY9DKRkKeLFiIZn2z6b9shEsXIqqlLY
crGcOGYDDkMnCRdqlvRB4xUiwj+X5N1rxI0vN628javhyb08c3SMA9+vZJVsTeAQ
lf5h4sT05Z2msZYeRXGCL4sjWdgUdHEKSGz7Q9feNgOtt2yK2IgQEitLjYIM5k8a
ygRwZIfvTdOzHsP8xFtLOh9OurzDZR71lFh5rXNOe5YChEP8FH/aikOJZk0DbkvT
8unxpFC0h7cwanpY/3BLVT/nEOlNiLBOM6d/p2jwzosZQ99doZrfla2eyyPu2BRe
ykfg7CC8iVWv9NogF/F7iTg2DniD3t4szval+gm49QNy9BPhfzNGpweI19sKf3Od
lKDFyGTmMT1Fr7hQfaUxUFWUXzL6FcFf2gVRoOU3Ycq435nszmDqDCgftr4enKyR
yyI++hd37k859dfIO1IYHyoiR7tDhU6p5vZeWU8VI1KLI67aWQ/cc5AwM9k2hHRc
hKn6chF3wjQq23E6V7yzQeUUPM+rI4VSx9A+uLYh/v/nyZjZepg6yGpNrHTFw6SF
VRmMHmRcYLNrQyfI1R6eUKAjBv/G/fxxiU6QwTEnF34H9DOsCgC+n13rtSvZ4spC
Ovq4vsmEXWxWbpB2gtHVAv9a1GNYMI+XcVPvkvvTZoCgbtNonW/S4p6PMREBs9AC
ocsCSvOXDGYsMaIs5VqgVsBxocUyqXL9kmUXFk6t5d/3GpGpGGYsPr+LwCBOA9cN
ceqPPM2s1jSIf0rDrd9+myn3l+gNqlxBaEsCXZz4sPsBbv4j5Ej/EgtoqF6b95lE
GchkToS1NaNjDBnMc9/Da7Z8LwG3xmgVgJWduRv+EQi2r/Uqcd1euPygwvl/2ahH
qZIjmfu/y1JSk857budXQ6RtWnogYSNKfuxG+qsmBrnDUH9aO4kjCH7OoDb6IaEm
M5BAbB9fFDMQaTfiFvDQPnms8sZTl0No972kk10IO3sy+lpxWQDxNXElekxMvE+D
ACjqwrPospbSz487kzl+cfb5EKInRapcNSu2TF3YqFFWODSviVC2s+tebSS3muDu
6okAMB+QtLBeDwjA3mHhQ63YtQsrtGbN9dF6m7FvPkWSFBgHv09uWgvC+5LPfiPF
fpKvBcBlNwsYmU9/cVxBJZXZ8kL9Ho5d3gMPcn2dxW9gtVNuYp+cIOEJ1O1MKlcu
idMPyU8I+QKJYACDaSg6YM+QUHQd7I8+59M4JF6slIb459KwvjJ/By0ASvvy8hZd
x1CVeVk431XOfAS9DwCc9/TLhTUm1q1GadnJ7duFNUKKN89pmHu1VCNx2L5hc1Lf
qs5YNi9vPO5Hl4no5FEfcTsmAYeiSRuuQUYGtxQWE20IBfISnPDMK18EfujRg8dt
CEzl1sk0hcriefnxjUtjMJKr0W+RC6SX2lDkBUSZUwVefmliTnU69t3Pigheh+Ry
UHaATkSuCfmkDL+F3FYF4Zz0nentRJyE8afFNW14NkKElgtpkNzbc9fPWZF3iMQo
WIxw2RAWNGkJ70qXSpCWWj3wI0dw4Mn6J2eQC3P7MvN5a3Y4ckKr/sfXlDUHLIj2
Wl2m190kYXTR7+/ziPNsqiJiwomKVJBDIQKLD/i7JZhWoKTmLcYeycQYVyMqiM7N
bOADpTtvvmXylmj76b5+CfrZej1620bOVyjM5lypQ6OBv3S+t0fc33tNcOsqxhIb
Gc68GHe7SEKH0btO9r6cVQRN3a8fdbnBp+4jwMqGZrBg+cqRT2DwxbRhN1kghjA6
Hvol0mNRCrctUiJWiz/vhEZpML29ctG1PWD0MDBlTeKa9f17JHoTGplv/akZpQTD
xzJssLfiX7RTz+iGn9RsOlWgzjZdRYhF3d3sA0sTwmnqCD1h5195yQS0UoHh0Ify
XDqkGaWhG+0ERmp36k9UpQ==
`pragma protect end_protected

`endif // `ifndef _VSL_AM_SV_


