//----------------------------------------------------------------------
/**
 * @file vf_axi_type.sv
 * @brief Defines VF AXI defined-type classes.
 */
/*
 * Copyright (C) 2007-2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_TYPE_SV_
`define _VF_AXI_TYPE_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
QCrj//IO213JR1mLxmUpDy+2odgtZw3C/S3E5vgsBkPMVutaOPowtZT1HlBujTla
K4mBdggOe4ExCN894IOih3h4efzDRbUcKt+g16RLPbl1rxMF0sp73qPRDyksj/Oq
/KxuIcgMIrvMgJjk7dlhjs1WAybU31J/KmsdwKwthmpTycXBo627xNUVk3u3OGmZ
gpTsyJV8Jzx/gzIZtlRIeZfkrbF14spbq1vt7yP1RqE9fMm9e6sBLW0xInkzXFei
YWvsdb9kBdbFq4xsPbAQK+HF5T7vifcpKIXzrXSQB4aRmQ46LBA5uvBbhQiTU/DV
1ARRa0bBtrd3V4zDnn4MKw==
`pragma protect data_block
N0yGuZm/aF7JY6NrZ+xLjxyf27eNLBFcRHqhRERFHJp62FshTGSHthJo7yC2lxpt
0+IpyJ3jPM+aBPSXqb2sDDgDQ4UUQkPSFsqi5gFgbV25PP6HEvfSxbZ77NimAvIh
4/RUGNwr8UcwZ1As8UFQ9N1FaUTQNxoN/c5xn4km+Ejsm/qnQayUIc3brfM6Ocsr
dL6TawKn0SQOHh6hkwfRIiprkKRW3j9Qri9QPamw0eJUNPb0qfv+tspqcFMMbns5
1JB9OqOTPj5pL8syTBX08xXpHHt5g+s0vI8oX7muRJo9qevPl+fgvu58J7JH4Gf2
gLorj5ZQ2AvgorczBZ3LNB1ssZiyBasyeW79SxTYuwCXY81MLQHFgdsovsxdUV3F
9J7f7JMbsAvrxQP7ub5exFScR31vOFokH84CnEnRVxUvl/fA4LOXCM2j4U/44IxL
JtYxE06LvB57zJOv2Ds+QtqZRbR/gp3mDBnn5sy1H+ii53UrlppbxincuktiM3xY
i6GEbPtKcO+UicNn7tvNChJ7Azyy7kuiyPzVfJ93EwHgQhzdxdw3br13EbXd7iob
hBBOTCHFRw5yAbK5D2ryuGw4YpdXEpm9ASv1sLjInBg041bE0IkHwtjDEvYgP0LF
lhPiCjBjS0B8oL6pFCbyXG2Au0kLIzr1PdPBAXiK5TJ+FXjP26b7HYen8sdlOkq/
sEHvC06pRc6/LrEsIGbRimKgiNbZlozj2PUfob9ph2GaEd5rh5PEA5cmcgtzEbjk
GvpAl//dvUewqFnAr5OAMAZMfeOjVXgU4a4j0M7QEAyWKGJzWi4jQIi4A1kRwdXP
Wqpw9UMtHry/H2K1fq2aQb/tXPP/8uKF96mqt51Fquo1CZPdcms/VMp95I/rcG63
wE5stDNN1jdd+TdWCXGe1BOn1HkNVmxWZ9SMSGgkBVJptFuD7RilKQ1GBH/IR8zu
6lgjqE9SYQyAHbARTPBabav18Wj+hTGxXcMYGFPcVFpYPCtPUEn01k6Irkgparfm
EZBuJ/dpeiKsdj+npl8pieQfkwlG1iWiM+RSFFwGQU0dVDP9NLV27OyuNh6qUwIz
kxeIE5K1D75TXcWvIybKKQihb8nw7u3nSHciDQR9+8nmzKEI1z41kio+y4FI2W84
Vzmy0kLWMUpLUw0glXELVQfVdVK1NpCuB0uxA2+UlDUdUkpH21hF1G/BIuopvdBS
Jn4fPdwigZpS4ZlSLdkWUQgaKHHoz/OpRvTVT/wmBxlod1PuzmoMMdrA1bimEnWG
bRFsFcd3hl72cALu6wogiWtrTDXtrS8P5y1rnGVkFnHwLMXLZuq9x9ZyTWsmPlAq
SGSdM5onEL8CKt4JqgIUkF2yfvllTzjE9aDCe6ntA1gg34Ta4ToGqF2/QTMkyLuT
xxr7Zhb6h3lLgTONVAIpDcI318vjRBeQsD0J+mz/e7Z0Tk+y4Jn+s/tchuVXh8CJ
G4Wa6q39p8oGyWvGEXQ/j23Iat3QzEdFyH3b1eub0BIQ+cGswv98vjkQBxQkTE44
C4Pi2seXuIcssnnXQBwudhOv26CUgIkVEm7woTvXl4kh+lxyOuDkZwGgrJD+R2c1
KXAtY5uZUBFA3E+JRGZnrOccH2yvySC1EfYxAL/k8saE0f/9z7Hx9nQQzdtyEoFt
DdmgWB//U8MhHvJln9M8Zsffyk+0bIGG4/Yj3GVJ0yZPetgSW70d5YW7aRHvJcvn
ORB+fP9YYlFn4Y+eYohFRqGroWe73E7dZ/b/ykfU7ZGx7xRwvUezHSHHMTgF8eFN
sSUWqv3toRGrTd6TcTrYKL6f63OOJ/TbWBEXtZjodx4ll7TsXIU5Sf2gxVtCLljY
JXpeFKryudFEMNL9DtXwjfVJiHEcvXGXGmNE7ycR0QsSveAmAWFqwjw7jpzNymMf
7pLKSytW38TPnT30gCoMAgdQfT/HIcquGSiFG7HqdGCSI+R0KCnp8+uycZ1zvDeE
/H5Qktol5W4gQOVlBczySplGA4Gt+YNJdP+vOYWbNt2oyiUZa2FTNZ0b+xHxXNuV
1LA+Mo+Dcr7uWdkX9g+i4pAEbRWvIlRS0CG9wguiHTuk+G149BW+ZQp+noZMDYlv
OIMOSdLKuOSduuEYqFfpknW4ZpjDpar+QATTdNrLIZddqwDTAjfOl3g+jsdLCdIK
bIJVe7X5OsWEETwdc/3SuTVyDoy6f/Vx/3OfMHZOm4b9jab/d85Ln1BwnS48l3WZ
CelnBT462d+Ga9MiDvFlv4Fj9Tx/f/3Z2U32KdgelHEZqTpYnl0uyhfoceXQccx+
egkXudHgI7D2WIYmc+8IkPC2buIPF2fRGhYN5Pi2RlvuaAqZeXpMED7RK+dehUs/
WSD6EO7KU4Y+O9Oxa60rDtlO1jXEnxCWF2LYR/xwAa3aZG3+vnPaJY4hXB8IR7Eu
m9bFItVugef3AsuXt3d4hpTCWFoc8gMcOUS9gp5ALxyIc8yXOUzp+0Qi4nYGupZT
/YZ8T6viOinCBMmcmJp/+bz+3AOj/HhiP5CjfWwr9gEsnJgNZ+cpt89AgzdGSzVN
3QPyNFeroONp5OOKjUqJ+tQCfYtFuvvHcRgxWtIeOo1VJYYCe0l5jWT9VCagZ7En
hKKMwjgk4XM8kvu0L9gdWwngLV0Zpkd52LeCtpcZ00v9lWDxZuW5RNrR19aDfQfJ
Mb4F4Hl4ppiopN7tGI3I5PygkD3TkKFXPCg7ZaveRtGNB1FtffhAT+1VcRJaMJWe
uLf/28IwAl4Vv1cuTrn9M6HZ7MgSLYCt3nGP8g3UzHM96i8v6/SuJvpGYTMStXgn
dpyt7NnpaQ/G0AUGJjxeSVonqOreriXRgavR1F3BKGKBR0kOyqJSEyBYeHjj/0DN
dpLfh/OUd6ajbd44bhF13QwQJtpDlkkjjmH8ngqo+lSkEQMpjclKeGor14UoDKfi
DV1Ag/YPa2ap2SZIySztweTMiZW1cCyjjyU83oKUXS7fC3mMX0Q+skVAYgj5h0ZP
itiKrkMOqTMg9ZKpCWu+cjE7RgDflTLacuKbRzEA6cBWYvUGtMtItBQzmmM0hwEK
+Ilt7pwAi7a21cXLeXNAxvBiUxaDVOTwm63SN+VRuxjKQRTclsNJb4QrLB0wy0jK
NHLskmvJSzK22l3FSzcE1YWBXOGQHcOtS7eKghG3gGlSf5YUXV7cSxkNPoEWB8oU
f8Wko4JkVnN8aUARmTFwlukZ3R2Qzgx9SM4rGavyrGawycq+qyhXiev2MykQ7smQ
dRfPlDVFAC7SYnCwtNYtUSIqmwFNudv/bTRmqbtHvOXKB8NV5eH2ZkRugOZA6h3H
VlHM2r/4l94K3JUGLbiBuK2jWSmuyjaKw+f474hnveyQUqLwEuongtwKzqm1zspa
5ORUPV7lk2HAnRHwkN2nM5th2e72EUYvjGMMKbsBbZGyx/iazaQrChLAD1PaFBco
+4wF0UyW/tnWtanRt/JDm8P/RUqjCcqWGvDxtqN6pIVN5BWsvyRnz923OhgJHKJC
83MdgZSJx7MjnDlyZLe0iavK9dBQ4fo69Vz6Zg4AYnMXEWeh5kSVNGhtFOfXQX4k
WZNGVC9XKIWw2uKeIiXX+HOSM2iGzhXJEJB25C2BJapaadLQznWddAMN22r5TB52
Bjh/jcBMPedc5+XnTxOB/Is38SiXaPCRLl08lmQ6kKpGgQgB9wtCYa/7iYJ5YOGP
M11JGvgNiXkoYapff2jjcDDd1ImsDZ84XMtdNE+QSHX+xrMUWAi0DGqkFsrQ6zR0
BqzI8M8wamCR5AEzG7lE3Ag6ZN5orSu8+bpCXEpaBxKGW/cR7YoRkErLxA1t6m5K
dRwReJJjaLw8Dd5hzD9by8WLCzKm/LvTKSy3IlepxK/+g/msH+0UpOMQuDjI5zGm
MokvHztTlPMIElh74XOOjpk8RwMuiENccro7ZiV/0pYSyWhBDVgrtSRGe+jrV9UA
Q1z+d+qbdi3VS38uaY6SipTWEb8UaKnXOG6ooYUwaV3e1gus7L+m6VFHI8QS4t0/
fH/kJTtWDFWqf59hfCtG896S+2FxBNZCaWpxxKfH5iIyG3iJR8zUaA6QbVThPAXs
iZqIKeKJagjPKuoseSb2BQUxdFfjOP6I1hQYeGRLO4B/ZC5v1allr4LqjGW/ee4e
aSXB1nZQNcSnY7mzETw0KaRfXZ5m+/qxIwKqIgHOGU4DQoxfHwEtrnD/cFdUOfeG
Jei+eQAnaPwhvBQYckBkcDIOubnH7R4h8K0gQ9ork9B5lPD0QHE91tBzmZi6777V
1mrjGrkQ4fX31wxByEj9tUUrHhol5+FjJG0mKIPYmlUvC5aw+2erI5blK73qd0as
0YLTR8RImtS3FZ+QDNrY5+re49OKgS+ta0KUn+xBqu3B/QBvi7xymLvRzNF7E5I7
KF0QN4b9MTFimKI3vGY+eYZ7EBFi/HWlItKe/gwQU2PZc5z4qe9Dt6P27aISWGRs
/fMiHEv1JdGXi0CgsRYbtxSo6hQ3PKg8pfG+y2NK0LkUqblNQHOE3UudrRHV6ByS
MUy+dzao32J4dj5j0aYXjRthzavUqZElLkrKQYVGt67AxJv360d0Rlg1HuI63RPl
L4ggkB2EO/b/FM7Hd4mLKTJUq2cXzP7hNimnMtEYXaIuomcyTpzRMcbDygasCpTn
YxpdIGtSaJ3fu1gXhnBseCAi9Juaj0KHwTzV0Plg0cPA3Hw/wuD8p80G3BEf7ZGI
MY22mbvrXmQSxYgjm4BHrtJoGblvVoLif2bdjg4OaSxptYEOAkGuqkeexL++cy+t
CDcpUeuqeI+o3Vv0BqcUujelst2q2GTlsvLA9GvOttwihq6xU4dtcQOjIr3AP24d
qYdJ8O/apyB9ftL2+y20fBCyPn2BLZDPxPNsrXTJBlQGj/bt4xGmQbnhiDittwt7
G0mb4ssP2GwqkVlB3b2kgfkcTJhKbD3UzBAbSemEkFpp/OZCfoU7PaOzzm8htqYm
qt8wrSaCY5bJo+NrR4t9pitUEe0g7YZhnA4GpmxegytTHjpbe2CzBuKdVXsNGh8H
aG2URoThzo6nRE9lXREK4H00eV23JLe0uVnxdUV6vqCpVqn1B7TtmrQovM2LFxS5
ZXGCYxmDTJSKKMqDl71plhOnpxvXwkLBjo5Pie1j13Lu2HotN3XweKLlzS8h2xmQ
Dax1D+ENTEs/s1T1RQ84Jw9RYtjVXq4kpoLx26v1wufZF+kHT9458JmCi/0t4LN4
Zsa5wGqnEvZln/b/+BGBaMWoPOCr7EeGhlu1GS1BUeHsyw3ivtny+VvA+N51CvXl
ajYy1EHCHhGxbb7v+J7dcpJ3T3Acnnt6IvC2J/bSSpLUMkRVa4j/BYMsjKCIRx3h
NkOmoarR425FGOm1SYzwoaxlDnTMWDdIWo9FkcELTs5IVWEXoTjihnFBtVri/0bS
5iFvSniGMXz8zv687iesHIwAf4LTNcawW1t4dCkkafqQvMYxaoujra4+Sad0C9pB
4PgrqLwx2uoYgeMODMhbV/PdhugD50CUUSxmUacWllb5wjAtvXOYNXjYcXLsKBAL
G7ZNno1ThWhNUQswOXr7cTxKQjohdjZnIyXnXAnMPrGwrv6sgzXEDQewFHmxk//p
dZJLenviz+XzEGf5eRP3WONN81S0g+TzWZFsXflJCJZBbr7iD2KuBLeaxZD+4yAa
Uqy8UxIVIce8veHVppnmRs6N3SzNAYobwQ8FTl3ZdHfQO2RMnapdPSjXeVHM3ApI
gRJ+5ir/E+fBhb9FIN7UG9NTeeZTPdPAH3FbmNMF7Ewsdcaz/IcVWKdwLL29MBf0
NQkctgS0tUxkJmMbHhApw7c8yTvZXZuNBh7kXLzRXxdqTDnCy0ob7/Gxps/P2SBK
fWYVooK8o1b7vnuoN8x6A9s1rpzHgLFR8+q82sfaG1jrYLA57ugX3/493/ZcnQlQ
2ckXXdaSWzu2NEC6bN6Z9YUtuZ5KeSMSK7h/Qz82CM/lOfx7EcjXj5r1K9uKl7Nd
Y1yhGnIwLcdLkZRODJZhhsn5FlOmaPzMPkgfDuG/7XwSyaHlyrzpr+27zcpfibEU
+P23HN7EJF0rwzBKhZQ1rxBBe5t7pxpyp9IKaOtQNkqXhfMXvTkhBVhVnVCmOMXY
mJgpXu1PrvfCfDda1xzE4xdOQiZ5GmyJmFUpmKIXDtZLxOeWlJuqrUtR0teNZp3n
jQUFiqR6Ab15PEm5Y647VoEhHSCaVEO21ZNzx4mg6wp9TUu4nk+i1DgN6+9s0H/b
/zV1Utl0V6Ul3DAO1sdGjZ+tUzqT/wGQNn1+frEqguNmDU9WGOADm5SKEVu0GuI6
4qZN7juef6qMPeVwrESAQ8MZflQc8nmoDbxRqY9kbFYgPjOrpY3h1mkR4y+OrNSg
Uh+rz57wiuZfZfRIPDmByKEUCFdr1LCnC+oEpac/kjJr2C2hE6UUNYgUCTIgmPgS
d7V9gqIvJt31+ClbHTHFWwofRH8F708/pK8UrNu6h3loKphfhS6jdGi1O9PFCQt1
7/A75ZniacJ83sRKmubODbWHNkHhdpyIti5hrrtDFMa3Ly0bSDaJirWWcdoKSNU7
KGLcA6QLwihDI1NbKWh0KQkhQF510IkavS12AiVIim4zgN2QKxzocaZG3ACssqx4
Atjh690X0MIXsGQssuRhuEyK9BVSZH6kXx7acd1C38dq2f4czE4lQK5uByrEFaxj
w2voGoeR75CCFxjbHoh+BZJnBDMpo10cTbRSlScBMvJE8qiS+jKlBKBvyUJ4Z0fx
JJ5Pi3nwn6pGkkIR9X//yT7GlUHWtLuaWsZ1zmfUgR5OLCwXYMiCF6XJADToG9is
Qg33LOEJjX0KbmuEWT/yaekLSNB+6Vg0tr5nbmxlg4OTkyZ6k38YJX2CBYpztO5X
45VtziP7LZZTQjA3+HHJ0qJyOMXWiawXRQo3LALWcbz+tZ2oAf/1wcKm5mBboWLV
NbHqEE6dsR3rsLxfGV81e+C44Vmx+UJxtl0D1010zXSdOP8ZacxRdRcdCXJ2r7EO
G00d2At2kBsAMyXoCzd5uYe9JdHTsgjIYT6twJ3nYZgNZ1N6NTZoOcJObxDB94dE
RLqLFCK/lKnpwG4PBA7A9I7CCOPCplwM8TXxrY3OxyA9+iC6N91pihHgeqpayJIn
yaTOU5RQIbK1AlwgAuBd4sWnfn6Ie2Xo/f1q83doT79ypchGyJqt0WrjF13inIyr
sNeCiqQIDaBM04bPlP4RO7kyEJxC0o76CPjb1W7jocmAy9ClQ1mgn+c4iPUE5gOr
ezl51P5Q2d04PIk/u0+WFZk6MBhU2yZBhWOl7N7rQYzMr/VmN2fDWZkq8zFQT5X3
fXBgnyFq7C1S47G3T3+9N8kfobP/eFmZGxgoUdgWxqu3EcJJr2ImcAcSV2ZUIlk2
gWXYe2aywqhmt7ESiOeGbZZAdKDj7WKQ5ir2p1VLUzKL0ixoZhZ6zmU7wkxlYq3p
Hh6ZEYZWqtNUbp6l9GtIgvo3UICxiNUpz0qDn26helEHkFQ0kva8u38YAIFFdEFA
Ih1DG5xvWGtz6BdsIwVyJw/E3x8Jk2YTSiEDkvc6pxgjNilXTZijdLcLHz3907p3
OhfYfaOaHe8x0lvVm8qENXwCZXxKdX28s45UXGe7HBgo8HFS18jmNlIEG73lngXd
CUSLvNyskblSiMYrU8kQpntk7iyFJeowFmcLv/NFQoQcdQ/AnY6H2THmcpL0MwSk
GLWuvr1hE4e1qq79kXU196GmxXnKUUc88q4SR73gls0vVziXG+ktOQeRKQpJbBbY
xDI0kFQPJ5PAn13cRS3W37ykuRmdgnGpj3qCwLaYM9nnuH6KsU3aB7L2mKPPZ+pA
/gRvEVysuekG017pf9PPL4ImgrNbUxxK0USf4/QR1+IB44jyVZFWfI0JFdHa87IZ
cU7vSjZ040gpSPZ+wF7sSmWXBOLUqLEQ7pJQmK6CD0JPKi5fedbDrs0dCeTwb8dx
IyJJjSakKtx1gajjVvwo01WnZeRhG2vQ8+kGwui4C9yYYCrSFhs1coRNIQIv+i4r
Ak8XDXpNFhr+h9FJcP1jc83njaZL0tMk5B5FuMjkczxXGIh/P9LOX7bQ4j4ahFfn
CQBSIPh6TLSdAKmZkyiEA+L6YTl/YAVL2RKHFzuXzbhrWrkGzysQoDWD2ohyyAeg
4WC601lY51OK1FHGBgJRdxyqehA1HzkdchsZ3D6iIVXYDYs3mh3aPGkvIJ16IDgP
v9WsnHi+fdBkvehT9vzgURqb0e5qJOlzA/Q264vf1JjU8EuaVTQh5TSxkAqk+4cX
XACEFxPamDvTFjB/jJW7okbVBxZ7CNqwwvxyTP9VWRJkcP8kpoTYcqUX8lbMiK2q
GsEe0PyFXktz8tcZ/sRHS8wbT28E3WZfrro3SEQ82zjFZQhCUjRLB7nlMyyqRy0f
A3/dJ/dQD1+9Um4pqsR+Pfup8hs6UWR6d2cpxPYiCx4xBHL0zRtGgQvGuJtiwHSI
hFaES8WqS+NzPpRn2cLMwv4u4WCUHaL3DxXqKt+Bz1kNeHd2dGH90O3hma0DzNjD
YL4C+JBJmbfkvcRpdwX15ciEX2AcIfBXQ6CjqxAruFe6X7f6kwwk6BD4Ke7Q3hML
/9zvY44OXvOs2GfPFAHrahVQo1UCMpkmJmaZ0S8T2tCtcrDV3nSsr5ZHhN4Z3gvf
Uz7I2CJjOL8+MX5yZ3Po/zfZ2jRByEMCvNcum77S1UU+dlbrShX4pEj5uIZGBO3V
eNRsScS/ZYP9Wv+xqDCt+5x23Iu7m4hIIapoUHtfDoHIWuhaIzhckCQyQ23kp0hR
TF3afYNx+PAbiJQpzZuZBq5YTR1VxHSs8KirwYwN3SNZ8ex87A5Kc7GbOjJjYOtn
UwUA90JlZgHDpM4vt2KrwtphqMYViCM+eOUa28qyszKo92qX5hqhPaIdZe4t6rsr
ZfprbzUvaArYAHqrTjfNRQH+dsFDlsjEexIqFQaZtYF4GotFlgmTx72edTjvR7xf
NIdmmThZq2CkpveMH4YRbr00Pu0PVqHIqiy3UJUsCRFHONb1DbeYQg3g025OPHN8
h23xTDYe6M8y6ipioVNIHtf5Gw4C+nJaUNf3BxnYWwzSNa55pASj7eZLR0KJmlXa
i90tK0QQd7AB4u7n0hHx+wiK5Q8qZ2oUNah03hhJe43UYl9/WmT/Ezu6m50hUEOH
9N4mPwikKih2FBdi6d4uMl+Y5boEEazPcl6KgmsVVy51U9RgZYavfw+sWF5OBv8S
sf2+inRx22/blOwXpKG0xSaid7mQKpbIp9Zvn8zv2Et+YU9l4reN92pgfDHokGTV
4z5HqKoN9afaIgqTzTXPDKMdgJxYr4Q+sdtUPU8nVKcpuotRA6kTZUwwzj2EcfAB
1uBE4yfPR0JwYO2lckaFcypaZm0VC9AgqFP2wyrabkIUXLmPOT0IKAbODKRyVfmj
JShFp+B/0yHOvDCgVVwKd2GjbxpJJSYvJzz0mCepdb1Ny/1hwj4qsfw3aG0SkH/x
ED63pcPSmxr4LR294vmcfFcMg6UISpQZDR2/zo++0++IQaFS78XoghUpwUkm03/O
1zNUJLd/rENxIVgEPvqLxg65Ba1y2p6yg+VX6Q+fbjwIA2HoqbERjlZC5rDVZMr+
JRAn6qMkBEht4WrqhKVPpPpwiW1SYkAfIsDqfC5F1GJ6Qeeu3zNb6PMRm81jdDiS
ZO83VNYQkJ3fOVT1aS/ihSvbq0BIcsgn7+v7oAGyf0Pz7UaJdhir05PcgTwpjYe9
aimoXrTUUwOIyQgBtADzXhBQTeLU7gECM/AXy1Gth/I9BKI9o07jB0qK3rL2ZrUX
fy9SpTeVLYCV533YCNJlaS3x6g07nezKptw5dbgUxJ6NxlZ2tj68HtDtlFYtBSOI
bIb7/hq/QC4P+T7/JWm8u+9Db20KWhNleoK6UvfJKsxXNqWKIYmpz6Ebsh/4E81I
Eh3csgczDgyhaWukfcC1wc5RqWPDQxIVx7yGeH33HWzSOBRL4GmcC904o+fV2FnJ
Rc1j4jAFGMjLBRw9wAIC7Cd/K4m4iEMxls5GmIZjHuaZH3yikWYSdyL7q7y/Brwo
ed8o0jROitaqV3irhianFSMv+i1b1bc/i+pR2MTrpTtRtghJww1fKS3hE4WTDemQ
0ty3uHcqeELOVVby5ZNOrW6QkUsEwTGVVjC3jqr5S8cfSI1fwoJqlyuWj5nOA1qL
VpoPO9F3nUq+QkTvOqNZu5TbQD8IUKpl/pDr2wIIu9AkphCkI/IDMa0U3Mrhq2vH
/AmVze1mUGTpOC9UHTZtnKX+77bM8B0osnbAtfoC3NZo0Kz7DNHUlANdMl26eZ5Y
og4TrsrH19Dqek6gmyLNaSevIhY3ieFlqLn/jQzXToot2U855ydEEyNZCSzy02Z7
8rWYCkodXClX4FIptjo+/rpuhjfWg34PYP2vKi6K9aDV/gaHDnTAE0LJ2VUkf1d5
S9Ch0lt5Y8glM1rgw6peNgC2JM3ldAFAQXtPV7Ob7qALuuT8NqzLceqYKsBdih8r
cE8+vtvehNVqG4gQJ9IMg1kJhVZ6QidSBynN63ySCAd08z9hfGtOoGGQHG+8SJwm
7l6jKZotD1e5Zm/qBhSHf3I+V5KJQCiWHmyiNL2WIHJnhXGTxW25hD96IzKF4Dak
f8mgrjtVU0BREXnKQmb8IlJzSZk+Dgin8SyJ3ydw2of5V1R8dO4MVA0IiJopcsFM
qb7Uetht3sSzDhWT0/xlLqgAldjYfvzgNUZVOlaHj5SmREkxYxb4JTQMxhtijYRt
VMPc9gY+0brGBosNc8N5h8vOyxwFCdHHPZx9zxsvYAazgzA7LcQuOUa07V6BAlQN
+id+/VTObb+q6ZHVqpXNKTv74f1qp3X6jXdmjHSS0Gtu8cgvZLj8gjzrwgemZppv
e/zdIOvX2orR/zhO2hZ2j6Tgy1KCXWz33pjJ9sLQGEfa6o+YTHhF3Yqu9ud1NVUl
h0jot8t6dE5gJtwPycIkfOzoO8hqH2sSzT+VpqHU83YEzzVcionw99x948236q9r
uLczbqVArx6/CLX0HsihrUyzHXsy5huSKGEQQ7nwpb/Z0LCgkrvGynZvXuo+duvb
g0yZRiaNabraZrAyQJdnCw8ZZnljtTjRrSTtEy2/tgVfzwDUc5YO1Iml61xVR5Sz
1deYiUmpwv/SFewpJQHEvWnYz31q7spbJHRTnz0SL8/EXx2pPdi/tnilhlgS5Qqc
LYrBGXpy8HW8dO068hsyKPhGo0Uavirxwc8626r33egdf14GM5oCZBH1Bl4PgY/O
1wDMlrwH2eqMqd6PwUj2Zw==
`pragma protect end_protected

`endif // `ifndef _VF_AXI_TYPE_SV_


