//----------------------------------------------------------------------
/**
 * @file vf_xact.sv
 * @brief Defines VF transaction base class.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_XACT_SV_
`define _VF_XACT_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
NALKS7Tq8aD7R3fnBhTjhZA0BYUzZ4OU5uOleRBGSu38oYTLb/kvgo7OtQkb3f2z
1id4G3TqGOxwwj09U9U44k+nj0sMnuYWUgI1YlQBCWTs9b92IuCI2VwmwkAF6WVv
Dpgw4IxA5B/4Nbzfr6XoK8/dueTOGpkdFeM5JDpsvXOvSFIWQuFlL6PmYXs8j+W1
UcTeRfyG5aEb0ppjc+mgK4+3rns3igPVUy1/DvO96BHGAgUR1sRhg4IKHUvfffeJ
5A6dHH6YWkKhKMOLX0iYiLZWpMvS/EEQ4en2Zhz/E88RDkNZhmZ3sySYB8VIpDDz
3KHO5+GCsV6cABfiDFYNYA==
`pragma protect data_block
jVWWSOqSduQ6VS9o/M7Zv9QU1WCVb0dB8NsqnTqP9VzsR/soVtkOZBYkTpvu/sIC
II0D5phIr1ERiDRbmW97rU8Oj1xyaqN1KyGGrN2e/mib+lzaSdEH5jYZfMA/f0hX
IF9u/1HONT2D+etEDUWpWSaXbFnsHZsdwUWICZcB5uzll6LMo0UIc97EjLTvSKxL
W8Pc3UHLDpv9mAMXgBaKTzRA6xRyKaVlCiOrPGw5PVm76BrC9xpbqGdwbE8Ts+3c
IKmLgIFDxFApOEfHh40oPFPG8yBriD1adchmyvWvdO+zz8EHP+4M7tWbu20kJkDj
kVuDj5CV40r2TABjtP7PaS5EDe7oBrvmeWL4BVGiQ2QajT9VLQ9bAj1eF+vG6UsK
2gsEP7sMep/LDxYlNWub9pnY+OVdoP7IgbUuRTUTfzZH+tKlWrS4ld8064zW0dXT
57p111CMjDCFb1uFHf9JZB/sBqvFUePoFlS0qaAfVA01IjpYUn5laXAhRu4kD9QH
5Zno4xje9zuTKiRT9Gt2Qw80B54WSTv7HMrIBOePTUm/IqzpD1pT/lWWplYAZOQ9
f+XH9+Ah1h8Y2227pXOdvS/3ZP8jSNOFjJwCi+o77FeirrSimwES/5dI77Sw5Rlb
RnmZGv+OC8lU0DXvNdSe2CxObcs5/bGnG64PhfVt2r4gQSuRA5nGjpF4RRlUz238
Z5w/znDrY+SA0/F96jJzZukxdr6hmJgifJz7+mo+LNBrzS0LpSEb1JmlFctSe+xy
wI+NWDmdBVEIngfVcxcR7UofSBPe4f/sGp5o1hwjQmjas0+Dgci6r6uJAgPhTs2e
wXa14bTEVTCwv1B5IaQ0wl7Ka1xZqvciyXd85N7jlkFfXjZhuPjTjtdYawti/Z2T
8fQOd9FqiablndRy8iZjXBjX+7/T4x1jNMeYoF85GvCo2l7lwRx1jK8prV5PRIgj
JWefAbfYIL3wmDav76FjMIEFeGX0f9SJ4ed6stBJJ++ee7spl5nIn5hEevTKLiaZ
RQYdx0NZv/WKNnoqciL95XuCAre26G6AFyiFl9SJpd9aD9KjqBTUAF64yRuHsOjX
pV3q5G4sLF9P+axvpoRRzg3CWCbKx7Jiq3fOgx3kDhnTs6dQKvIKSdYC1DRa4idu
uTzMKHwK0mfqRjbAY1/IYDDeZmyOgGc4bBNVrKJHOwJDp9U+7kf7YtWHElFOcwdj
XmHwNnGQJYTS+x3d7N1JMVZ+AdLRRRThOct+QE5Hr7cKtj+7ErH4jBX9soYn4Aii
ELyJ82TFm/S47o54x3k03+nI1e3nO8TJ0Cxg4OVo10vcfr/rchk3wFMLAfCo93l1
1XdctB5ZENrEMjv53N5P2alHVLPs9FBLSl46HJ7+Ya2pOz8tINj3cdiySOiuDOOO
9urRBzAokiP1fg5rUWYlI4Vfa89hZMC7UzboOXunXX92GvSXHYgqH3sXEP0E9/JO
wxchwcg0O1dHlKGu/Pil53UlFDuginMXpwymlfKUc05+dyDJ7gdPmnwnOn1YfZSx
7oOuTdM075PBb6IGW7g42WNEUduMSbEiCl2SO5yeeCnkZeoCSCe2l2eCoL5pK/JK
x1tcmy+D2T/zUcrqcdPlFehUJf9PoA9Jfg0PlWZIfGsgrB40LizT7bMYPf51fDb0
eaOjSV1QBqJC+ygJmoD3bQvRz0VHeKrFPY/p+5hFcfBBQKlW0L9aAFySCMwQNB+F
uhKcq3zaFwZJsuvHUCrfZG/brizYpy4sB/CphoBM68uFwRA5p6aWb3n0RQ7RqaeT
pacrWuNx+mNeAKdiL9yPMUSh1DXR5J8FTfInPEQ3QLEE3ikGXMK7dd9S0P2GGfAz
FXB67Zafiady75kLqNsf/uB7dsQXMOFDaDnmR5CzUKBQJYAMyDDXsF6DIdPbSBq7
VunPGHkwlrAVkqfAa3Ox9zaB3LzYwG29HuOpawrkkp1QDgLdV0anBJswlA6bmmxR
GPxB7SvQ3cQPdcZXVUoXu39JOcXaW+sCNw8ODSFoHsFdRK/erY6DZg35ee8uVvIn
DFb1f4+jo5SJAnBkON8IQP9fYHz6ySexO49YlEprlHAuyghW10OUI+LMKsnyJAia
gu5Uu0GTlJfRJy1MNuJCeyMCBq2FKoLjppyXN/ja4QQXf3JcEUdHUjcn0+n1cX01
OPROKTGkXr1MvPj7+W8o1U3qhBXa5ME8U6qpJWr/mN6JMQdrHHyIuMa5n1XT0zZu
unF3lj0RDq1+ylvwGhxw+s8Jq+v6pUSv5N9gI6cXhNfTVwyRuK29aeWBpcR1BGFR
xBbVz2Hcf0+PUWJjNPqeGA8OkqC2kuH991uerM/jmYtjy/EkQwAly0Rh188c6Fnc
TKXHG/L5vcwuWGN7CtuIcAl1kra3KPXTIzCercBSRtpRCPTuV9rHV7UG32D7BZa9
eTfC7+58lqRonF8/26KMMDe46O8gKiCuObVnDAkk51gi3I7On6ALkchdEiGqlHUq
235fM42oS4yJXgCBPQCibaRbZVWk/AHbJ9Odob6UEghSkqyOfZ5j1Wo2q7SeA3QQ
ldpbaSLqIv2/NGIEO6tMI4yWehpxh/CNJdiSSk1u7olaww03+FZJWxd7J9O11XNl
6TOLjej7bkxxK9BCK4XePk/bJhcSqnqIzBs7ezjeZsSQZwvAf0R1On1O4FGQa4bN
3Ubm7Qky794ATX5lI+llJhrKDJlhbBk/3RyBhRAPVFpVcaNAYe/fF/mL7q/EZIrw
+xOdyQuJxxqWpBnUPxPpbwvYFcpHHw0M9C6fO13zS6bi53Gekd4jqQ/edZ+XB4ye
NWgsnk9gfe1QP5Cdq8eD+lNnnBQuEjXHOyO+YACLZjgpNvIEzfzhQA0jVAHizJSB
EkGQSYkxjfovdZpMT+WElgd0DL6skdLVeoxs8/x91u5cFUhWIh6eiQjVVMgrAIBN
1NS1PixNvevPIBSKglg5rK33MXyEzPvqDoqZZBuywq7IIDpbKoSSQF1vD7AnB2ca
JuKUxxhvgNXTkQnWmrvEtRP9IUQtAQ5c/SqQmXQ82sYdPlLa6rpI7F69gMCh7mNd
/PMf+4a7SF7m1WrOs6Jfjf0eY9MO+FQ9HD1TJKCFwaqF8hDrQyd5ptEqIdXXS9jh
aSJAVQkdnLgGSD/l8FcW9fleVhTutC/pjjTNkCfjdTBFzekW1kKfgYZgDaQbMcgn
W5pjJG0FAia2KflB6RVPUN+TOObQWU6jU5ruQiZAIcaGnXe3N2/yh6UsSSYW+I5I
a7obNakQ2ATjy4cgHxBgwhoVPaswfknWu207PPWxvKORrObfY3MJX2VviX0yO8RB
6Vcu+4fyGSXpGm47r9fjG8y1x4rVLynwhSQzGP9HqYkAxvAKKUYyzLiU0GIDgvB0
a32+F6U6Q5PKNkjDg2E7OUtKDXV1cGMn7/RzA7Lq9GQzOE0d8MLAlYEXwyIbN2V7
TANrnwfMD1wrsMUhV0/F7Zz72AV8SSIXYzJK9atKrM9g6add20LDxTRh1bVzdcLn
hAWMeaQ20e08m3C00gntfWSMQcmRAVc2GJdpV4jRWLOTNp9HjAka4pxdHCB2tYWd
d1o2agA9HEmm2235FtZktb01RTt+nMAOEBQ+dqNECtxIFpQPfi1qXoWk4kRbDp0Q
r0VHJ/R0Mx7pCM8qaQsK9mtajfL6LS96WNlkd0AtwHZO0ww8jJX0voak9gieabpe
BUyLB3pMYo37FzBp9cbKF09/yzeWMO/X8/rqU7j9vZCaOPXecP3i1YaNJ6wnkA7r
UnQ2INd1Vv0kEqUi3QVWLCiz8lpjTn6MzGd5mPkKYzikw4RVbgEZC+6jTgZ5t5dj
pwusTGgTl+D8We+ZQ9d2O0/DWaJLTl4JybyYQA7rT7CFkjhwE5aYJ77sWEilO8uK
0wpum8D1X+Gh5D2d4FlIsHvTcBgLuIJ/E6IkGlSs4/RxcGzxvl8gkQwkq0l005aL
2J2ha9FSb/Kjwl8VHJVFGuS00WKmYtGYkbl5jRhedEV2ffLR3oVUoHjnQHqBPo+2
/pIkYwAHeJmPOY66xOPt/oq6Hi9ToJkrTKXdTRhrIYd9wfXAVHB2xiojt/RiHSiu
zOAeAVPT7kPBXvaQ8gn1XB9NQtymY7epnYY7MqCFx6xX0En9hxt9aexGXzF3oTxN
sacs3xGg4ZoFeElsDbLcnPjylQjCRMBThT/KQuj+pJO3csURmxPjqz8PFEbgyE4w
f6Fx1y/IA/Iq7hrPXT5e1XND4RVSQ+uzIB3npPMJ4i3oA/NJ6n+LpB13Rcb4Y6J6
RqXT5zcH6BQOIv0deOggzFKOSTdgn/xsHgCDwr2nl0u6eiaRYoCz2El9L4TuVPUX
P4N2DtdulsptiH3+WWLmRCB5VGocRe9t+r9J9tNX78aLzOP65u1L8OVrxJCDdwY2
Wn2F9GGRD9igfkN5ZLFGGzmb/Y9j6/wXeq/RrkrzFX+tkuxfOtCA6SN+Pg7l/dW6
QIGxKupIH7/Qh+5i3HTd6snDzR/JqGIgSZ7Z5lde1dTqULh/39PQ7gUcqwDhYvj0
kHsLEo6E8z7yOBczZ2yoduPWM48azTPV9Z8OS/77K5DuCnm/6nkDr4gAOYJg1wME
WXCrdauc4OKPNpmd5O4VmCeVVCGA5pWT7VQvdtVcRpAgJKT5IqH8jcU7DgB9K7OW
7PImIjfY2Oc+/3kG6jJb5qsDxh+wVZEm6yEn8qn/+5VpOQ8ZvYU57Ul3CDaxWQ5L
gE4DBZiYZZ5U5xiyCmyb6PbDd5PJLkzI8lKkcAEcPwI6GEaYBIFw3BMFUdURAsVm
Q4sfAwK+As8pr/Q4zW4SqnSftoSd2U1KN6L4UiaBXUgILSFHQZklUeTOq4IJU40G
oarGq5qsbXrVsRspKl+zI3sD2pqxXvgY5mdEP3JbxyTdFCI03JGPKgVm/pM5mhWg
4Cm36rufgzT6jS/1FlB+e+Ztj0X0cBXrV1eNivjp2vmjXT3QJnfyLJefLxmHHlRh
DQZxOUb5g4WMNpG1SnpdH9w5cY+5/FIxq3lAGf/fFwT1S0H4DpkQH/vQ8jnTFoMc
5AnQ1ZQV/AveB6z/JodffEHYviRRRW3NEQSEKAMlEKwE/5laBqZs15ZhqO2zDLW2
HkGmY8Q+53B+tXZF88BC3JPiK2sOEkqyjUPzLBZdcQcH2l8kWd2LkhKOGgFQaULS
LY1B6fKoMV0h8HoWzCJHz2tGAVwtN3ZPJ8FpZ/8qb8mB9yQbnkTuElKAgeNNol1t
8Wx7Jme+2sfygR3e07e24TdNFqc7g0U7fKjwONMOMcgIJMsFqsa80JzXbP3uJY4E
4E4gz1bjAaMY1ELvZgugZ3begGz7+Weja8RdZOdotA6OgNMVqLhbbj6nBpdwx1Wb
hNtSTOR5vNyk02rSnQKupKjZ+8/2m5e5/eC0hH0uJY/tYLFqCdenpXThAvEQfDuh
VPs8rY22CRLkxtGZGmyxLlVqhjmv8o3UbSATBAIzW5NFVNJuASxcYxaycaufxpU6
sI9ZQzKmewrXMCfeClu4dwViBdrXyMwi/sKWGSEwpIrgOJxt96W/6VbsRbpcMThv
YWzSA9NpAfVbYJZQycSl4WRl7o4Zb1jUJ0DjeOY1XLHFNaVBe1aCQ6v8A5P1Dn3U
Emxl18bB2V2aWDqHGH7Wiq5zDvB+G7eh1zKKexOn//mC+a+QHV1Ms/3eiq3N+2D1
JKMf8CbOj/cPvIVDiJfSqa/Z3SOSiosLHOGNfT12O62dZUO2eZdzVwBETLAoJ1Co
kVnxtm/8z03DkYW0lpt99opBbRofdI52TJTWbEdulxOTUEn8epd+FUPh07liiWlQ
Pcl2+GKlE+bukunrEuxpIuBexNNbg6lB9o75ylIyjWqH7YqsUdKPcqEfrW1Kh0mU
vBr5nNaE5xm3XPyFILBlWMjnyC6yrIras6jU3n+NvnSWAwY7iDPJOO8OnKjMK43u
4qxN/As/Kd6dhjm58SYv9sDbip4sVKMjsX/GXUcpBmYy6DU1Z+uRJDH7kmERw3/j
LKJZmnXbVI3FPm52Yok0oaaCBhZDlJdgVgfuBnXE7voM19z7Hb+wrPKEZVchaGrj
1nZ+QDzvSVRD5fnnotjmgktHmCtp3ceHTQ0k3FKOxGJgOZq4duC0SsMztPRfTRu4
e3hkX4JMnYbssmcLUVJVlVxsZe032hXd5W/5KK33bsqwXC2aFLpmLO1SDg8Gy2d3
0RetHt9eQS5TM6NeNYDQhK1AK9fhYkrZGCW7yEIVWWpgV/vHMoOUAYOWaDwAw3Zx
wzWylMms4FWAeCRq/axmot50LPRz0mE9MjjortroDl+vLJQyq4d281VO7O63XpKb
JnCBqfHgBctp0jitlPOoGLRGX+gk1B8E5jEF3MsnJhu7anvXIPzVg+kWzp9L4j5c
lm9zrbB5tBbjLrhvyJsieYgmWEFHpTGdPXfABUi02T7kyK9o65EHxlKSFKH6mL34
rF4OhJaZQ9tgsiCVLTrCISm7ni+n1t7014ZJ3IOu0s/S5q81R6QKRfJf3RbouUg4
kxoDQgHi0Laeq60Rm9xClFn9VWJzvBIqpePf85CIWjCEW5ObACqRVm5JkHaVEaMa
5y68G4O4PWwmlDjh2CZag/CrdT8BEjLLVph+NN9aLE3dSi7+SlhD7cURsK0Hm2/a
vXLPXyy+iWjUeu+mqRLpqkWteG6tAuna1sD5Dnq9fdWt7yQy2utNUYgkxcWe/Rxg
wurDNKXXAjotUojRTAfEO6GjUvQzSXaZUvysbChoLY1BQWHwitInbTpYhAeGdwcs
y8wTHRwAX1MS0IsXwuarZqyYMxhtA5FHk7xEguEJhVKVVvowmolWzFU45TLIJO51
NmkQdYk2XcETR3K6dmlM7IlLw781rOpsjwS/cQNRW67GsHjkUGHZr8QD8nvuBdfv
HlNE5Jhu1nNXiCy0SNWnr4wG3GO4OARZxlSfkPafRLfmkzprDJgtqPvoscfEM9fM
cmvvy8ueBYCJUIOfzOcNJZqjk5VD06We9izFsPj93f9fH6sZgfQK31Iuft1Sy11H
LDZnqTDLmQJofayj4oeNOJwcIh6gaVcDcAAyDx5vtM6SLQOQllo3OvfQQp1ZliC1
20Ys8s9mSdJDZ0TVUXY2OPDz3MJFbaltxCEDSWeJu/0qJA91JOw0RwL4KX8LEhr5
aS4Ptai4I36nC6xNQcn1/GQC06qHnbUyjbQ30GWeP6H5PaqVmcaluG9Ev0Ixxe/i
iVgKrljT1sjgIYHcr3/K5DFkZTfEgRJNOoEc3qexo2KsrpyovSQkj7otJ0RG03yS
hooDlcqF4davPcLRDIcr6bKjmKQei/r3O8ptyA9Tm+F3RTepA2Ckd//bTxXj0yKR
zAQAcSDAkoGde3YzfhwXGmX8RUHadh+txwPHOVnx6QS2TZxzcVIoeXbuwABWo6DS
f4/3/LGHGbtXDrIxCsKz07zlqGNEr3Kt3ZvSKqiX3fvvNatnXQbnUeIDQSWfYnCL
Hnf5Sq6hwbvg1Cwx4ILW/nV7nduXdk9EHldQk8hJ7qX7Hr/nARRBI5Y+pwpSBhOl
+BRaY7yEuFC2x5RJdhzwNKCviKI8SaSdxxfQPIe7IzzmWxwDTzE2yGTUbI0mfpR6
X0Xjzslvxr4WGniOMWivLLsx6x1+mncmT2o4xZ4zI1/i6ylOl7lBmP/Waehchi0Z
OTVyYdsxdULdQgKKS414h02dG0YRcG+lPGSzYzog02Pgky0CyOYjX6mh6rGzNk8G
lD56E49q9qn7OsM1Ecwl23uxeTcFDuTd0Mo6VGWtPzbm48vj/UFhMC/s6uUjqG0P
bHp6RXquUnx+VKC/IGj8NETofLUglNgH2MX19Ng7VcEKq896VE8coPYANQ8XEAr9
yjUzgbv2LY8SoAMsUOqGgjdzEzxrzKNVJdjQORMARM+aWvGOaoK7BPZVmRmkN9N0
z1a9ubvKTE71fAcsRuw4yifWqhhoMrq1WoYPT6PuWzKw+w8pf/juH8nZaSNHQ3Qb
wFQ1RcHqX41lqKlM8un25z5YmSGpgnIop9v2Fhp6XdqQ3NmmMbl/kveXQkQB/tV3
BICquv1G1+pIHrfFx+bYYJ0h6w7SLK3iSmWYdOpv/+jktUqsNH0H/nArPp6eNses
pa9df/ZTOZo/SxRr/eVXOo9afCVUgxyaMDm5G6UGdwNsJCFtN7nT/b+y1Nkr+Nd7
7QQByneIq4CXl3e10VXGaFFWUmYtB3PbXGL9ND7Pv5dxoyLronhDBCHUqY/TR37M
LTyVXB1cTDDH3dd1sSmciuOfrHvRWDcBV4riCS6L2SFQ2JCvODgGUI/Ox7dN/gLr
PNTSs4s+WmF+d64dWAij7FB8PVKYsrHwCl4g4yZpyYAbHIqOzoPLdkAzwL8YRA22
mJEwU4LHmgQUKe1wlh5TN0RPrDgFBCUTrgS5iRe3FvaHHfUSJ5CSy3gKAqqynTwp
cAvVOKMnPyMH9b9I4jqkViKIDZL8xCKLmRkxmnOEhaiBbaW9cop1VrQimEx/BQ23
xMYnFZOl8gHoGdLtvf45f+dhiCaq5kcJ4Xw1UHUbtJw8y0bZfYzXdt3eRoSnVYU+
VPlp98mBwroNVRpDJHjb83vmFVtJilW0MTXfHMBsX1P9EH8HaMx5lOXTUKByNZb7
Se8Oja/qIr+rZM/bNGgDIwl6gOaIg1O4g/Pik8eYS5xzhw4mrJ4uz/0/x/3E8aZR
fXzVb1RTGXliuishsE79/GB0FGzXeV99HQajnqdFQzsERJt3ZcU82i2F9i5Bu5lg
b7JaycKsOGtgMZkYHc/miWQoi7mUXOq41Xb0mbjAOIw/r/XFNqJ1thUhh/biOgJY
3smiTAoz8/Sx8G4fPohW+xbrKblSMRY3Ldrp5NB8exfbfXPHCuMx51cjQ1cJMPEQ
ixPeXcFeZ1e0MUoRK13G9AJ2bAxZgvxYj1mR45XcNWv+vydYXrUqb9f6B6rtNIYv
DurYYGeVyirGpl3hNmGsHGPbQVqCMC4eQRI9O03hE/k1UfF3dOPA4lDwOY7zUCbJ
r7n4RhVCyCDNrvG009tif1EYD8uKeHuPZvRnFgUu/6+hWTJ+31zd23J/Y2TDZ4Yn
vY3g8dwhbD3zKxgskbTS7ggd9h9QxOCvf5hL4VVXKUt+/sDN002UJ7sK9Krwn4ie
Y6XNr5wwAXPW25HdrpnSegV9KOd6ngmc8zzJoIMjsJAcssR4v1TaeyJQaPlhbA02
uWc0bG8jN5C29dSpN3zE1wDgd3ZN/VVQEGnONvvRJhAt0o0ZInIiJNNIufo2WA/8
JWoui2463zSsbhgtagoiJumCqNEGfQLp5xvsBv5k+Eu1BfQZf4LB+8kQr2yNXNZ2
WZ2r3Y38A8k0Z040RRqKul/w3Qr/++tEThVWR87VZ76fr1KiLt0MHzmn/uNzsdWF
PbCkRk2xYoZ+0bxc1+3xPe7xSZoJgdSWRARDbvqPbBrddBa4mNKHAk6RQ/F8utR3
sH2a8uMTep2FyysRRTS1ZvpjZYg2NalUls3H5iQbHMtb9+NnFGnvA5/uhZLwJR2k
YXndaZpPgGk1soVa3Dbchjzo2wCgS5o8a2wTgW9uQbJbwnVSUIZ8TOIkbsTFDSoX
1qLkAPlN1bpLxuHJBGKb1H19t9XGmt/K0hggWAcWIjoPpFjImp/flPGjCl4U766n
c2STssLhukGeIXcZYTWQInKnw5ZhP2sPT3KNU+JJnFcfh56FkRIPT/3FtOGxPVOs
SQqLN14TWH2A5xqz5e8GEdlwtMCq5B/3N1UAv+br/NUiY8mSMn2rOh4MWekd6yBv
1srvUq1l4XAZgx6sDnEUTVKxvInzT1HLNYippF3UNypinoyvDX5wz+CCK/IcAPlv
sTQXjMRG3uX+3lE6OtW6i40YjJVTNJpHiIzy/upO/oz09C/q57vCXM5hmQX8nQqk
vKudjsXR1hKTiKr7nGkTRtZf56eRAEhkCUZ7DScJGDdWjZ1cVU8QIjy1Hdu3hUxd
/ul7M+UKhrzqtIGvQn7nID1sNOFEcHbArFFmB1O0meLIzQa35cYJbDf5FUdFlLMH
V6i7koxpCJFNh2eKB1FrYmVjq9igm1e+8aTGV6aBVO6VLCvvx7+5tLh4+4USUkUX
HnW5ivJaeO+w3BXR+pMBitVHEDzinIcL7mbRnN7CdJ9dnO47c3Kr+NNOpSaXt1z3
QgajVNUkIQdQF52ejdOLTm/4csk7OA/zr+faO9u9Pl6sCcD/7w2tbWjvn2Ejk/IP
LRB+l1A2X7ePYgl2l1qSMnlyy7jWJ/aagNWyVOOMDtlr2Hf++w+Fi0VfIiAT8QYR
Uu7QiRvYEqcLvK+zDeaOIrCS5/2TAu4k1exqEFBquiyU5A2X+JcMvrywVgVnE/ll
TAHiTwV6Tc2dQnhjcfg0dmFzE2Pn5J3qyQfpv2tkV3FtFIZbyhCkyedirvvXg5RF
EaukDXfwqREel4LDomKu7vWlREStxpUQkutz4HjDFyu5mv/i+2rSektTX1sHSFpg
n1gdjSaCx02k0vbAJmkNVguRFM3ivaMyjaKzHX4jiNXb3ako8e5LrRsns0l3QCLv
IsZowYPg624e1gC2EUrPS/bemMQFTT33P3n9aH6Sc7wYw/P2uzUtflq7kd/WowhH
+f5yYUs9k8ELxiDJL7MC+9KTa05XN0QZXpV9b9F46LunIUCQMyWODh7bjm1S3YBY
gMnGC+ZbM5H779NY80YiHFVDvSjAq9Oq8JG3vDh6jZX53+y91LbuE9tK+il5ZW4e
aCPbtWIyn2T7k5Bn5kUK4lqt4gc8Y68eJqSHTqaHXHmud1qa0tGDnR2P/g8xeqSo
HNVB7AQHUSV3c6h5zdwpLaT9pmO5WT23Vw9QwgwXC+xs8PxuknmGicbFFmRnUsNI
7lLWm1bNlcOTAW/LF+bj9torPbt2mnxhXpA4cfcKXHOpheQivl6s2ffMUJOVaQXf
YCdmoqmVyJ6DjjtJLl/b9BnJp6/DkMFjTlLLjX2dYJkvR9rmNN0/WGIo0xQ7XT0V
PmcNxrBl9d5zYkBqqbBLq3D94SMHCIGlkJ28iddm1VuHO3PbPQ/21+q0ad6EZ+RZ
NaZIAsaJTbiiDORezdWxuPrCW4gReMfbdDYtTPhxOwNpaeKEQg+rUHihWD1jfyKD
R1rgV4SNyYZ7q8o7Q4QEuepzZ7LEjujg+PqBTTOfKIgemnBybqSObARbJgdIBxE2
g5TWhXa7ZTwoKyo8ZE21TqYeUptPhOs/wk2U7o49yBh33qtJZUPzVrRbhPPmsahg
zJeSyu3v5iy3yuEkqlS7OsE4JYwe1eKP/nsDOKBX69qrrBYKDcciIjFFQkK9zdyK
WqY999O0Bvjq0PCklVN+GYVMkbYh0wiz0gUpDub5P/h4vnnJaYDueT3OhsObcvGH
ynD7orFgal7qK4rADrtRdyoa3HulF2PZPyHt4vjr2bNeEeGmy4qakwoUvuD5Ya3R
XIio5Hkk+3abhPo3adwbi4CU2+4124X7YjpZnnmUI5DL5FYKuxnHA5tJwfiTbca3
YCHlNdT+0tQoQ97rclw2vyHtSAYtIrt2xczmlc349912l0bKhFslFsKUartGeEuP
oBiL9fAmmqazjpAMWaG+VW1dTSKB3PJfAo1ETEqCzfNwPo2qs42HevegIgxtT1Q1
pXht2eZjb4tsULF2dv7FbeUboHkq3urNSi3bXl4vjP8YuXohNnImMwiEwIwiDq+8
v01EPrQy6/Ch+urUjEJKcBlB5GRQ6psOnljQVGadzvSPdr4yFiec0T0PcvfxMCzc
8oaRgd69+K6OZIo6yqEZ5COnoc9Pg0ZF9RYbe8bmHw8FJOW0+5jWk22uBvnebIIm
u65b2LzcEcIqR3yPd299mo6+55RoIyXGQkBDwlLq0navRdrbhlg/iAHRThKmMrFK
ZRA5dZIEXiRoOBjk2GtU9hv3+ziQhT0DuWxecybO2MwJcv/B0MD8oJo/HF/AaqEg
xw3ICdtxsBffMj5knRgYd/Ox4YgDuTtUiPlK7B4j+ulqerLxopV9tm3Ot88mSm65
S2X76cc/6Ih+GRYaYfsWar4vKG/OB/TcewyueLf/iHZRevfdWCta1NE8bba8L1hy
AG2z6XzcUShYnkiP9LuqPKhlXILPNju1ImwsGp8QbVFHKIubVPDKavMnMpeQDcky
YkzmwGx3Gsto5vDLSR7RCZ8PImlQ9azMgSC/UsjBxDZlcAGoqV1QVr3gnkJ72t5v
cBnrbXczj2i4nbRAwmp7rGw2uv/V9uTkZogn9aAyQzhnneQwYdlXWPf0vXpY8GKF
xTQedw6Lib/OiuK0S2R+tN8tUJNN6TPMedJC5Jkcohj/211ugWQcWxcDS5ZDmtNG
rXIlL1SmfyJOrCfbTeHbwMtkDVMg1KLLNdS5G1FL3oc7l/YX6dOmUpniC4uzQhnP
mrhtyH6cNVv20iKe6d5wynNLsCJnTYNpBWq1pd2PKStvA7HT2i39uiviLE+yyiS3
ChnMIi+ZgWb9rlCGvmH/4DjOInH4Q74NDONKIWKNi/OST5sp/djwm7/GL1c8TFG6
3vlIOfia0YKaLDKgzeQo9xdimIwb7322k7NLjTvdLe7TLqIPj0zlfLOVFxqWPcFt
RVYyRrq7EVPYSCHxfUa5UQ5Jk0oHpnV64rgQbZwpPAjCIiDlegg8pYknJJXFk+zF
QkOqE427qUapHrNkbfkyNs1Dbxs76AUEhCecttdbHIwdJZ1KeHbi7gokOig+vQW3
WOjE7Wf8yf/XRQFttIRz2tJDawxaV7n7hAdpos1tPljUshceeV3q53oG4eZieQOT
Jmd3mFwJ8YS2rmt6pKtXftFiGZX+/D3E6ZXDjMhaR8oRqrPQFtI33IT+MMiqN2Gf
73mdJnrBnc+SARm8pOb7qU5ozJk9VDs2kkY0szWBGhBfU1giEwKb6Tvwb16Cj5YV
9ds2cMJW0Ezb8TukKvTUm7WHFpIb5W99Cr825MZE7L1zNbVE/DfuYOIczIbCD/Hn
5s/48J59/g4ifZ4GxLBwMHjCfu6hX+KUm302wOimFdzRNBIFGZabimxgwxhmPSqc
aVD0AuPrwvc2bpMVPyQGhDDQRDAZ5m8JPYnitZiIe4vstERsY0+ASfOjBNFwRoBN
riDo1RMxfIxX8uaKMAHr4Y3ir2eXAxrKKFhjKFrOv5goPPcPWDRu2cjGPIaK3vtf
hRYu5WwIvKsuNcmlrh5uPVL8hn6xU4aodH8RXA47qcpY851pRUx5c9KnZrHvIfEU
GrbyrN+tY85PvSpihJPTJnXg8o+pLjChC1YVfXLVAstTVCDrM5MKZdcyqQgbhyla
OzeF8doHpNNFIAta4gmQtdGw2QZTYNTTq/+cNnMzAVx/EdlqfBXegwLTh1e2/4nU
Fa6ceEJ4Usdry99wsbvVXf7krZpD0nDX6EC7goYO3OADiFsvJ5QgdngOtVDJs3DA
WBy4EJlqI3u8yhAJBGp0ImArNWjI3gZY40cfhelv4oWdK2tzhWetypqYlERKM4V4
Ct0RMHdOb1knaY0fmD0zftXDG1k15sT9SV/qTfNwr3x5+oqV0a0SvBcoAt+IbMeX
fnggvU+5kafFhAEjoNcRjDDdokRR27zro3GwcnwCUMrpoj7dZtOPjMdOoWJlIX9D
ZlIKIRdOe7tE4wiI3/1Gyi1vM6sEisiFQzKNodtxWVDsIq4ag1ohifmvQiaX/0ks
kmqAmTQ52PHrIXPx6OaDbrYW4YU4HHBq5bxrKCYRvQt95iMw0MrtZO5UkKV0F7Jo
syBLDlpJEcaDdNebscKLP6da9ETfb0rOq96QlYIJurSdZclOegSrJ+/3yoN+x1DN
NQKvsAKPaAR5ySZFB2gjFTFj9py8x2TbAawW7ApXMGUkcLHAIXbKXublWa+iw0Pi
BkLeGpnWMYZ1F7wyONBSHE/vy9UDd7FZFdwZhdtg82qaEZOJcghfCnNMrIE1UNNs
Aax1GupSdo3uhuRz7Pe9y9QqRsOsI0iCoKlpsvBsiGAHoqGVTY7IrUX5btf1jl58
2L1V+Ilzv6g4fupZoEtbn5N0XDMgE3csZbnMC7hiZ2vz3hKFm1xSsIRPFv6SAZMo
/NdJoVN2b5JAUk+wq3Jr7yW5x71zIiZaOlfH3XsxBjwLjgLEYul7jKwyHv55KgyB
GsCRxZGXJMY3zfS/DE+HfpipFuulrC2iwnn8IkevyNOmxdhLLXSVwro+oMVPN898
fJFIxI8KCNveege5JgFdjHCU6BUsRJKFiKBgyRs2+QDSBmcLKVYWm1TvhDXB/a1T
gkS+jDMakgBRTCHp5yZ3tmEwcMdDPFGcTRkSSVzknV9x0+i2rDbMvtqr+Rfvr5/2
Br/wxOy9KI83OhXjCgxDkToOB/I11TWGT5bVbK2lMximfUn+OBtsPi23xN/2s4ww
7fB11lVePqSjnDf2ADHqSwXwdafCmkYIWIyoOVxq+zGQSkauyUizTnwAZuBffnBQ
rWmISkx84EPG0xzSN+AlVlZcYIujCYzVBiaT+IZUR7rgpgRnRD3F81A1KWBH5bWd
Qeuln+RFxEBpGwJ8Azm83E+IZUf8xoTu/47mMN294monVF5MejzWwhbPZAOqc+vW
DGdeoRqP4MA0NJxu/OgATGXp3amNPLHrUR36AYJJK56PX/LWSf2xSPzwGzbzjHFS
pEZ8YwdgdJasw//NM6zmtxPXLmxZpwUo0QWLSltQwEBZ3S4QF2DK9HehZW1LweHi
TigzslrA2JGw0XRLnDPvOYMNgYJm7vMyJjNnlzPxnizTO1v1hCzQ7rQbnMg8Mitz
8EsjhAsBJgoSwvhPRsHgYl0zKjmiPdx27hHiWlj7EQ4eO0GOQFTBqWrhkAcmxDR5
RUSEmm3kLjC9/YlY6no/4PIlaK0UUOtv7EoFO3DDZABZyzuY/ZXdcBHE2T6A0SBk
Gh/AmWAutqJlifK31/PF/Pv35K8fUKhlMYbKDTLPFLLzzYtE0mxf98RgQ7tO12lx
qTQ6UgKCj6lG5txYbkqymC2p0q8+Ys2LrYsnryBhi9iWdGCkvcociynWIZa7updC
Cbi1kKSljz8w28i7ozXI9XQDPrGGfEP24uUNgtODPVJCIbllK5e9Z7ft4snOlLqf
+a/02S+je23gjkg9bXM3N5ybSwTegY/qmMbi/et9tJ81MWxgNriM9G/6LVt/pXyI
k6N+ZLkcex3EC1hbDroI3U51CWiH6TfUC8ywfmRFG2Tn1MB7n3cqlTyMKy3vg2fa
ubs3TrPVrP709IemSxyxekxZXfKUyAKxJfqhHASXM9B+0513qBxogpkTUcjuYR03
TyOmludZD+4iDJWfgbzpHBO5OFx8MV8WdjM/Vmmt9/1vFvP5R6QyBkAWMMQcI5TO
WRvQgV1iEADrbfXqOn4DbmFqaxgI7AbehpdZ6F+GKVbgGWOA5nzwNNeTS5y1U6Up
58zGvY0lvH85HdF5snbR+9IuSHqU2s5ZO+w2Rl2LM7IqCJiR2tzvL+pD+sRzWxpI
5xzWZbcV75yuOaxe/prlZhV7K8HIoVvWaNbUZ57ruLLyVqWIerKPTc/rTViM1pdo
OWqYEQaOcykcXl0ftx0pTv+soJ4wezh9Q0c2sdCPTO0FX3muEy6AeJUjI8jBd9Us
TKf0h0VTYQ+Og+DwpM6TRxL9Vzb29/rYQgkcsC1SX0YC/6sqUb5LsZrktxShHEmo
8j/i3fbCjnvwFCS3/OihupcSjakGjgvrsfTxK1QPIN++UDM1fOOAVGIJ1SH/Fl0i
y5jr35BqJWI/yVzCCKt6DrpXL9k17VNd+lYGKHZNQco2y90r/k8kF5geXsIW2au5
zOGcaq+iHeSE0hBjGfR5IiyHKpBLbeFiMwMaUcoG3vRShL9oITaZbLP0hvenMQLf
6c5Ae/qZO+h0u268nPOTLI2d1Dwdk2C2zAqjDIwRUTxMObKAX2hykYh0bjMEXWkT
bn7EuVKrDIX5w7ZTO9GWI4wYe2KLcMW/68W4pvik/WoU35g8Epyf9KXcd79Q7t74
tiQ6aK6OoR9YeQyRBOKgAHycxzjkfvzVORMradsCZ8Skc3qTAzhDZ9zgX6POVIU1
cGI+dBDbXZn0+I636KUQGR0zAVlL30k9F87XZskFMlBTw6HXTOSfbmc13I+7CXRm
CwNT0T1eQXNy5lyYG3c0mv1UyNXM1DT/gzA/NAkwS+8Kzgn7LvdjJTqBkLICINPH
XhC0pNtSd8RhNhY6ihG9EA7aNQcBbjjmH5zhp08cZYHYuXJ0Epvl4jsIIXQTUcsC
6hVkwzKk/shl0YC7kx4o/JKlBZIVQaXK/FmRMeUd/lJKel9G/cbp38wmZ1dLRIhX
aVh7DVI4oPCIbSJsXpNEPsNfBCU0GDCDMEs8Wgu7o3+NBhJH9TBbw5aXdtTwR3+l
++Y7JMp16Ka3WNgTrK1YAANwNvRBTBNkW6z4gDv8DoAnx+cY9tuFLnofZZE4Booz
GELGqwMBDB6J5tO6ADuteMzuHZ0R98Vu2JUeMtnnEBJ92Nx1Zgrp0UqjDyJwn+tn
Gg+JzYoupE6/a1kiTYbUSe9ZyP+8nmX8IVCftstOUht3rJYRaGtsT+iua217k/gL
8KCzLhoR4I65qDnzZo7f7PXycbVUo9KgeLo2F2V5pLopZhQfl1KLHfYRQW78LttO
lQyb/7G87OTERdDvvxuYBJvLHcTNMYmIhRL937yhN4OFOg1hqVBn8bMJmN4h/XBI
R8sgw17duR5SXYaHJ2Z5nk/0j/WZImhlsX/HE5z4mGtqN5yaPUxWUc3nltRmMjXV
rmmYuQFNmfuOhWhOYpv566EPGWCNCWglIrYLDq4ZUa7zb9UawVLNnG4mkwezbBwf
kqf5l6xZFoB9BjDuUR4Dn+DFvqwbbSibfy3fXTqMLbabvkCRJxp84r0SiBURTly2
hvWjqrvX3Lab27K/TGOm7kseezD2uu1OrrUnFxeydR08BjiYWfuCP/JLhAK+zsYZ
vIRGRd32ulLqMOBXv5VvgqQMYKivDWG4QGT+q42js/hmLM+TxZDqqHHmTm/bJv7T
HYZHTpcjhgNXw1mOLAjKZfkJfX+C4JRs90RwbMCzrt0LweXy+wf3jVw14QdCb/Xi
6BaJuqjth8H9XEvxQcq/1bmMR0pUdDMkay8/SSh0ClgwHT4+8knMDF7X+OIQUoNN
QHSxGhmlxzaMB8IJ1S6nUhBREoIjaMeN8NyJhTwrkUd4DL0CAT4gIDTnCQub9W/I
gBoKJbzTfjP6bi8ykxlfM4QeBgjLf5zJuV/YDAXpY3tOAPaYjcjFu5Hzd5ShIOOO
jfskz66VsXm9vgLh9iBbCMHiHlazAWmTV87CJ4E77EZo9VFPNhKhGW0clY1+wKmS
85oypjt9z46Euhb07vd8aGCK9btl1ISLzRkK8IqC9w5Mj/RfewMoj9wpCOA8tuSd
vpFXhbKweGrf9X8XDadGFm7lgTSi3YbNaYDRKaI5nBzXE/b6Z1lBCWWvDLMoAfC0
tswnwsYA6BV2VojUIFfOqOg8HR3eD4fPg83xVUeIC4ZR3Wao8iyJNJzrHZppUyEw
daY6JDhnXYhm80bLsyNvm3PiexZWCsJdjApwB2V9jljrEe6ic2u0XZ5PMTtTe1KM
8p2i7XcoiohiqoGm7LoSBR1PAHQn4yaIVsKg9IAAL9xfNvBsrQp2/tcTjIh8rkqk
qfHwqnM3/Bj4q6p80a2UjPfzGJuoh/PlPOJ72h4lE5TQscug622vORQClJFsKnlp
W5G1CYrjy2Q5InAMvhhYaRHdhC8WXGhGxhWViYabzYqxO9W/h1dHINGkup93iVDw
3nZpCxE5tLQtmuQCUu82Xx1yaNCh2TUHkWNSOIjal7CnJ1Co62FcLtyVU7wdowJi
P26TgzllZcw3etxuIM8yX77OMVYwUHaKtdLmBkSn9XBtjqgPIBZm913XoW+MI5PV
7Gh1GvGG3uhLWGCBlvzXH4wrEw66KzHQ0hvI1RMRhRx+QoXp1NGbUCGzb+x3wgjc
fg4PxVLTtF+Vdm+Ay6z6/aAYRSeq/zHLmbui5VyARZwwFZIghbRGOUeiiFU+1bEp
vkAjYiiebfQv4ic+hPzEnLvkY9lpSzrgH3+O3xkZ35o05gIUZ00Yqz4SqGGyeL4W
sHxSwRjfKe1CofXpNDlmdZgwM9sVy74qJvjCZ1lq7LlVWL/AtDJqADb2+pZSM40B
eKogxujrcpns+9ohsrvigrcSgVK34xPDcAgiKQREVcMC+h7Vetne2pDBeTOcIFcH
99DZ0DpH5kkvNqiirZETE6511KRDAgNigmh04o43s1J6bb6Yt19efdhUQKk7xfBZ
I0rASUbkNFA44LE24RdN7s6hMnRdZfgkQq4dLiRUGXLtNNH/1fhzs1icohs8O4ef
dSv1YNtJDTKDDW25CBtpANnihQyqnXrMGX/6TXuhbypyU/JnT9o9Xj8Oc3SOdqrI
LBtLuGN41Aa6oxgAu17a3wbE+wn4wqsCvFQ5R0yhguf0G4aMm82RKDGns/3ojWQW
r6rg0ma9YKgAWTSbGPmCBM8+4aaJpn45TfdegYohjFIO7wxnSFeTwz8Yw6fRmIP8
yx/K0plG7tqtQAITKaJY4QB9LAGmJj7fr4m02gzmwqJSyQXYHzq5rzOZE7+DZ4Ct
dqLRu9WVzRllR7FxrypCoQ/At7rn4cLhtcckRt2NG2/YXh7Nyytqktoobu5yWyCo
ZaULZ3wSqQWqH2aKoVrlGk6H1OMJ0mBBiPmCg/4o7UYHkWjJGzmGSnbQgwsJW8nh
n61wWspUj0xlOWiDrZgN8cct1+nEGOs7aGRoFhcsuPMYfxCOrw3rYWgsX9Zd8qPD
7RKqrRh8NEzQxZ9zapB/DgAMTcmo3ZIKXsNyF0RVE504UjhZBFn+1w61mYQpn6H5
dj39vZ95EXja52am72+SPaTtcTAHUvcgY9OR71Wd8/8v7MXfuD3W0sCEBs+JNnqc
t3+FLGZx55AzoGEfZmsENazgAwaSXqBUv0NfYawRqtDeBeY6GT0pnXRPyguXtA9i
iLgD9wUslILSudAXmBw7ol7sZ/OjpiKD4siQv9CxJOhybPAXeJ4dnJTvTMIphpOE
P8Zj7EFAWd6ntj+2lm1viHt9tBeaE95KvuO/6Q2izNrg9tEfHr/8ris5RB6J9j9V
SlXbe3WCONZ+SRthIpuXA3LIzMxWBVT+TCIyreO0YlnAjSdlF87SHZ9WvG69eST5
6vv6EB3emRm/w71OHDWnyR0a+KLQR1CjtW63jDVaQTXkHamGwZZ2+0pAIKWFbdaz
p4FSwwF/qGQ1rYH0k7T49gJ2Smt0G9AZcziX0IKOTcJ7aI4l3wlU1uSi1Ddasbkt
6vmp1w5sLqo9Tc4BkKmh8sBsvWH6hWYWzzcMneiXBN3mpNtfEbyFXanuT1/ifF8m
Q9dI028qalSjP3C8vR3kSos8OEasCJ86wvPS75LG9EN6dkUsag/Kc363qZvTyZqU
IHuUiEXAO20WaVCnMjJe6QMyLXJVYpZWwmot1D7ETJbWHkFmdG9RfaXQxho1jqbR
NWoIrrB5EkyAEBOJ/FCDf8xO/SWpOeQLA2c5oz1ndxHX4BcX5n9j5Ct6C4EK7Bqn
bWOxE6Rke+44Jw8X/PBsTVu3ywY0ozCKj5p9cnMv4l43ZLl3lIKV+ZmORhuO8sj1
/EHLuwTh/HUpZJv2xFrrNAAvGHC50I7j6oizHMVOBsa6NMyRoLa7HBHMTlT7gw+k
tLKUjCbQgeaSh+KG2TaBQhgSs+SO0DCMbwww2OOz0YoPxR6d6dRg1mVPkuY6A4pE
xO4sjxKdKA7us4GDJylGliPhg8aAMuILAwuRzS3hr7u8QqDTIlpZR5K+BdrJ2V/d
8B3KMMJV8Z8Y89AYChHXKScVDF4K2QBbtriTm0nc2q7lvZ92fcwAkGWj/+5kRHNA
U3EKz82TQ5r9Ka5tYCvWO2CFz/MZwwNSJ+1URY/pgN6ey8b/aFGLxNW2L9BpRz4w
K9ClyarTMIdazzQPw65PoLejVYDMqTz9bjiUQqZ23VKhX1Yygq78eyW4u2+u3oXJ
rXAd+XFm0G/pK51Ris1OUaEBfbyVXfPwNOqaqxHtq4dNlHuNqRvc40S2fSfE6Bfy
Xbqx6iNfyd3W7eGlr8BDsEhhI1g0S9DdkT5O+GvIlwDbIqJpLyyZY+B0KciHV4pc
8W9nAp4xzpWJv3gnYx/ZY8uWzrybbTGZTMfd3UHJ2JJU75WZL0rB0KDS8yLsxox4
6JJT0/lIetjYyZQomaWvL+zppHAFukcyywzSVQrKRrvP6109ooU46mQAKIbNJkCy
1J5EpizkuDBaTzrflWE2nSVTN336HLGwqm5k5ewdLffFy3sJMs50yOVr5Fntk/av
WBa2HnKyZStAqRJh6Uilyi1wz1m8bTilqJ6xDoOAhpoYyJbySsOOiDsYkyMvaz6w
B3ehMFxQ1NDpsHjRuJg015KWsxLcliF0letATsEf3AD1g3hA0D1ET14kGxotaMM5
k8d/nx82qyLVoO1GzqfaCTl/YJ1XDJ/Wf5Du9UYDiuwrLiQgTN2tBpqRM3+53Ds3
/dR3qskCOl4+Ij11Fxms9Ag9hgrnzjIzZj2xnXaFj0h7h+1nIYju2hS1BCiX07di
hTSFgYqa4hlmUEnMnEVaXSvqHiXlus3NSvx00MJ+CkjgtSorKjbqW4Q7Y4k6BmAP
c8g7l5Ivw2brHYXztZbwxsXQ3WNoURNH0mjhzMVo0v80fA9S4XQo6mDhx3Mj4zga
eTYwvN0/vz6SekhYS9dswXj/1pnUTqgIhVmNGS9nOvdUHtmIRpyHYMsYB5eO+k8D
/Lgd6Asg1VSnHHsRct0EFmIXgH/Pi7urF7dF6Oq23/YDq5s4T4oFF8Mw4oNQmOGT
mxSiwhjWjRtKTqDYiX+QXiYp4QzR8sE58LLHURab8e0M6A9ETTBQtu3pb2JnNpoP
M2aHRLudjkVa6j5U1xA5rWwp20bNSF1f0JDkS/e5xlvedgW7jr012skJrq77qPpZ
lIQwu9PncvdEwwmW2YYj7gnHDNoCUB0EgXZb1wp2ZQ6XmnvRxxuYzO1hhtchPV6B
wnpeO+SBxfN+N+4/03hNtHTA5tLrAEHEmueT52CF9uS1ku4lEB6zCCMaC0BVhXCx
1YE/4wmnZC33fAoCObOV24Oi/aGuXEMFn3pcbkJrhxixGp79z+4Zkc8j57JbBMAZ
HG/CZYMHVtUDH/mLCWpHxjOlYKzDmso4p+uF24MlZmbFg8MGFbTfV62Pd4ABC6ba
uUyGNZhOIdAgMi+p4CpA1yLN8tTUI4Be+rglQMaDq6Bnlk43RNHhWpWJHBtlU18O
wLmeV86h/1lMyQ7ez3OVoa0Eeo1a39PVn0bSmqLnxwCXWINXLq9qYnSjt04DrggV
6qkf02KMErF9HtwQ5ouw5UMT1WBMiqWOtC8eXjg3CO+QF+xP0A9cnHNVQmBZvSL9
FVwwzg7K9tCnHf7LMyXUR+YqUVUbGX0uGPu3eCvfph5DP60mEfXLYB8kdlYNaqMp
4V/myeCMTkEzz3yk+UPvKGdySvFuMmVm5WH15xACg5OBALV44QUkP1a3DQjcl4bb
Gaa1dq7weuGnmhq9ZFkpDoEqsrTr8jo4CMje1CH8tyBQ0dkDZYYiLaWpdouT3fxo
yGJwJgzAQi2HLhv3PMH7FSZ8iz2f1eqX/WXbNXSSakjUDLPJiAxXT/8b+KFpqJsE
VJqVx5ekaAGNgmM3rgYEWdcpXGb2HsPHYpX0T3oVkJEvp8HgkvWFtHBS6Bd4P50C
Crwkj4Qsj4bpmI3r4i3KuYnnuPh9NIADyKHSxv2LmGLi7plbSM/VTzTV4jbSaOnM
FLfjefIDYuHis7VwlgMFHaXySflH+rKRgXhgSJ9S1d1VmRaYx1eECZtRpP2/5t6+
YBtx198u/VSJW5ceQRC+IDYxQ8zFZzvVuEPGSe5mMUORus/PFjq6Pao38N7cZu3J
jIvwzkrMSI4B2dlotRVTScAtXGq5YbF6ttVq6jZjmPJWZTYwCKgddtgDS9uu/kmF
TwIQXYHpWhHnaUyvIKc3QpLn0YH2G+q+WiHSXyFNMlTvdNluQ+NqwmxiYlgVJIQ4
YQ9v0QZbS3nEjd4RNymBCFPIZ9TUVNd9C57azJaBdniXItQgqC9/cyWiR6FeYvwI
rNwJQfXdAzKOm6gBUQT5OojmI/Hk8vOrIvLnyZQMNtJ7C3UYEYn2NNGj28gnYZmo
wAoMOZ11LoAqt6ZLbdWWEo2rTMIeDm8EfFzV9zNmF7+iGwEUXM9Jn7M4GxpUZq5y
UTTY6vT7Bycy4SDdLO8p8/To0kLf6CnwbS/jbkogz4fSA1BC1cGK/z63gjaodCXv
p1oF2YgL4awfjVjSekDWwWZWVuRrZjJ7PbF5FTKaQVD2X0QKm9myFuAGa4xuEGn6
MzIiQxNTboVqoSUgaXkgzAhwIZ4Q+25nDHhsnqgAY6dh8HIoW2Ipbew5xi/naF+v
MO32LX11WucLTHTkdOR2r586v/+okSKjnXIdP8/69uxPrKw7uKqnVeVXeFk+Gz9S
QW0xPFtxv5N4Nfe/I8/U5jGD7MpMRF5tb54lpdEfLLJrbpFwx195Df+wr0B3XOJ4
XOsr00aDBsfMcquWaSMt5pLSRFzxUjeWj7+b2KEPtJZ6+L3+FBFOUpBt+FNE4N2b
RpprbkLJQGlIvFWsW4RLYSnlDxgKQZEmK5Vr9rkSLyF7B4WV6Xm9nhFAkZaalhsx
hvoOTZzmVpK/iEgbij28Jn0CFA+VnL6sKBgxUULDSqCMrEnhOslZT24dJ6o023ci
nxSFnzdczFP6B68JF8jI8x2e+qnwoOrN/rgwQ2EuF40ti1Rh9HLFiIyPdCzSNL1a
vxUca7gY34pkvDFwXa4vNeL6iRDUEpxpEr9WeFjpb64ORQJNM4VvR8iD1IxMbcwV
yIZhjyU02kl+SyuOokeV5O09f7RzPteSi0rPMJk4e8uVUCfIW+yTp39fQFhY+08+
xWEcwkCuK3d7nlKDNkCV+/ZSNx14EzbjhdgBjGL3ng+0r+6BccT6hdsWVOzyOo8N
xFrQBXif7WiNGXiMzAsuS+XHq/CbsfH1BTSOhzPZlQsWUpJQAUViEomCZBKvcEyL
VAN4IP23a1Z6KDnuEMkWLIb2epyLA2hjBQYGLjKGWosoV3r6jQ7vbk2Fcp/dwF2e
6tHKiZoyLxVS/l37DtWQT9mT6ZpG00piBtxvVjjLqsJ56755RD9V9UCAooOLTl/s
uBFd1ljwcsQ9jYFM7+oh3jwILsKUxWJJB0s2zY0X30Ypyk3U95282gmnh4AjGZ93
yURk8/RYrIT0+HQiwGJzAhTMPlWMMtHZNQUGkRdLOWjaCQxolnGlPX909NIC5Dvs
NIsM02RYH3ZMc/rKeGUO53gKmSbVdODC6MRbg3Z9koC7QnDKnDH1uGTTO6j3A/Ld
Hq4b8nDAIzGXUmMilgiT89n0SW2deeXP0aykYcOI+l6TslUecQVc+cT3ind6eUR3
Zx9jPcsfmKlPBD8KbD2L1Th+UixRkqvjDOyzNArHYGLjNevvRvJ+2CSWF9T9Wm6m
6Wvm03BlxdO/V/f/peSRdadqMADlsFNkJT5SFbtAs7IdLCoVrpoEuTKypjU0AJnj
chfzoMIak9Uh2LS7LFm4Wxvrn5saOcIC/IH7D5FaPF81dbGSNwxwL8mbjD9HjN2q
m5qzxumMcEp7JJrJFI/Waws/dkZ59lnFeFVEfqqrsrKaPx6MDT92Ee7RIF/kqbHe
kaOQ6jZLH55gxFHxWQmwxDHtV6oSkU+bdsYDV2uR74Ie8Qm36PaTdwalip/VAWsB
2MYasQgatSlye+6DZy+8M9fNFM9WefumSvZLE2bcVGmqsd7PJEVea+hJLHOYPdHY
beprpCKKS2kqgCI72ol0R2XEGmYaxWVj0o2NvpMCHq+Dv4Xv9FrjEOFHmRytkx4w
UzBPsBroPRufPWRjWaIASzA4tnFjDXoBMlE4hjWEtUoZBGQ2pmeIGE5nOiYbLdce
AepV2jwH0KisSwiGNAGn1Y7aeBCkb29gvzRJ11oZHy1qmQcnBeCGyksjfGSMmbw8
dprf7IYiYYKCZleGi01pdpeoFGvdOmL2mS+HomsnQ/VH1wevmk5KFUxlUPwc6o1L
EhGhCCda1OGSvNlG0OHRDbQcC9s8OZTOV17tFK5B+gAP4Gk0ky5NiZjQTomxw/aG
hfbcHGQ2hn3LFlzlhgaz9W4L+uapQvJROdj0gUq0WvoEJ+45UQhOxxpkHp7kbQ8D
T1FwBUPCg+rplldgWlLhorSQ/c0P5pjmccENWuBQnTJ+olbA/CwrATIS/g3IFnIJ
sxEOcQEGU1XfnQt/Gx2eMfWR1ZXE7MzCzrRwSNcU1xI8v61v9VpM0iW48PYK67Rl
+TdxVmyhPcDpapzO3o931TXrBhNGC0vz2QXHCRk5NYG10S/Ij+0/BjBC+ansKRPM
bdUCK+x+hm5UrpSO7sFV/3y0tfWPxF+0/QzVBFzlNjJYrtvNMIiJq4L1xCc82dXH
ZygeMobMcO5i5DCH78MsE1H5KXYaaNHB+bdWvhBzvQ+EBqo1YXEEKyEE2lLlHunC
+BSWycduJOUOLYgJ7lEdOQEmzBRRae7jGl5iTwZk/fEoMkERQcNz2Xemc9uoNlu+
YUeIV+oQp+DcfE8O3jpZEX7O2/+F5fNp0Ua8GVzoEySBnUwOlusn3Hu12xom0icD
dPoeAtuMuC47ZxzklxWjToGxbVqr4lgYGsLzcsBx3FPn+S6d53Z39GDSbWs0MC0A
LxMkgI8KsluyudP1yv8pz0smNF2nGy3I+18fQnaJfW8ryGtigv2WgW2muFQIuNzy
ZNKO9CSDm95D2JJXMRWAvN06D9S49VxcA97St2B7wPyIGBqPPDVTlUFEcyQyKKMN
MbD6LOBZLDvlRuE9M/StkrAnPMSwuXNKUwALEpXXIGpVytP1yMk99k7nUU7phQyI
DCtQ/XHAKVcSQoikyxF+uFOpL/mjAGU97YC3VrZvS+kamEEZnGmA+UC2AB5Ly/54
h/Yi9TPFMh1mj9cYfDvRuWQ+eO98+kjaZ+DnJSoeW4haWopn8cS3KXe0mQb0q1Zr
gRsADfDGdhW9cJwvzCpsICTEnw7Vg+M9qHZo1IYC8yYK1ZZ9l81ESq87sHXYlxLS
gQLMuQAyg9eTkePkUkV7837ynkEuWJTqO3wtFh6n8y7TgaH6MyuNqYdwoi3yv+5+
ny6SllnSEo9ILdOkijHOQZzvtflJekGZoV7+3UzrVZt8qdumAflb7NoNhACb/X93
Nb8JqtAcQWvm86K28YnaH7x5anAaC2ECpjtOG4rLq/IrFDG3cFbHkLCTwcyy6cL7
/3xUNUZZ/blPihizojL4xHf60H/YYS4cq+KvziLZb53pNw/PKvgaCDbrffhLDrCi
/VOX2yS2tIxkUpymyfbWvFA7tysBllYZVmztHXPRg+/ohEqag0NJkxgjrmuNvhIk
V3sJBTXyGVfTY10DmsZZ/uhZAffFThqFpWNsoXQzO71uRIk7gRejiqAlh0KSTNJu
rz9q5NYOs+YcnWD/5I3TcDokwS+XyE6Qdpjj9YRVUTXxuHsetRaIyiN8bBaeZqwj
HfgzQI/QyDxlnmlxCY5UCx4k0G2ARFfqQDONT08WHdRb36/0QxemjePDVzdrk7gI
Yf3SNuaQq5VyCRdyKDsX7Q0148QkRoVsNgnBmL1Ul1rDgNa0RiEl93HD4OxEXo8t
Cw8BFxnYCkwZ2/VWkx5abVGtYwcG+1S9f6EUDQ1kGNvFSV21RjKwCBFnlUrSqPR5
fqrfcTS/aBBKZ+1hiigmvg9Q19QJEufMSuZ3glMfpmpn2YI0rle46UrV1CPtqks5
jTl9wHegRWzReQDwri675RtwjqlPsQPt/1s4jyeb7GpnQyEKlMIkgNjwqJW+AWje
TQkl0U8ModaPUHejU9sOOxoajrRFR2pgR8eyisr5KeuToHscakhy522qBihjrnee
a+EDtuweCX00O1fJk4BV66ewqla0xyRlQ7vRM/so8i3SMcFoL9m1sNMUX55AmTsD
fGTc7XczPGGzYgGQSI6N/yq8/vtk73GqHLa9EDzyRzN1FLn96UhoBxQr4Ix1g8pB
w7eKT8k+BsVDt+WFtBdfV6mOZrjFaagtrLcB0TCkmr3xslmQtkJZ4z0TCI79El0Q
STtzAbdNxK3Qx0L/oOMoZAfSKruKfQoHiapek2hoewp39ER/wJuBlaPEVo+09bmY
Hh9nxMc+9cclWvdz+bchwXUynao6/1zX+uEQDSe3n8+pLU6zd6Q890LvR5DIKRZ6
GfP9wVwLszrIcCnto71wO0ghrTwNBVEQOhoydzw8De8OKeqphZHua36f/FmLbv6w
DkaVdQwoCMahOIv9sFaph6VkWpYDguzJO6RXbUdjtJ+cgIFVxcijzcYWuEFSFMu7
4xrRv0xIjjaWKqly2hJJpQQA4ciX669pkAWn4q0Qf2RTXsbkZPRhF0LGiUrT1Dvw
QpMOGOpH2VztUQfMzxunHnSLeN6Lz4xJGoSQa5Hs6Tio+5ia/bVTH4vIVZJpfYkq
pAxxDGQS6uTw3sZ7D+ezD9PkddVJTgog11bVtUVSbjOJ37tksE6yvD0uziE0BQw5
V4344r/V3ni3yucTjjGt1Itf3D21/TPXYBx96d0D3YlHrlS5BFHfbeBaW6zHhoug
gUSkebkfQ/wxqTmyMHk69/5YifkaugljWhPWU8sY8SRmr3oOQvgUHhmhslUO2UGh
RlaEYwfC0oeKyM7sCAYjecoO0NKika+dWCzW5xpfb6i/9/1mjfgUOlur+5HMWEKJ
0uibrdLHKb3RPUbAq9wTyhbBNKvNYyDxb5S/nP1hQub+tGVp4fFTdOy2EnvbWGYZ
kiibiT+vf8dutaeT7e4MFtZ8o8dG/M2M069zyBVQ7G5nB8ZAAdLt9rtMfap4pSJZ
W68FB/JaCQSv4vzxVGMbJt4TEwLjqDLdEyTKY9tb7OpabzWe0LLTvGegp7r4l/sO
lhr3+GdJdpf8/v/jNgD0npJlRWomSdZd5XWIVab2yW7jG+TuFFTpfbiCHAEkk6Vt
xQBat7bnGH3hizG6mNq7eHkGsiT/EB1NrPfltAFVljiA+RWE3JGNzO70odZb5QXq
VRLDyQ/rkeYCO5BVjTd8j3DeVXxEr+83q6Bk6yGFuysrlh/ilr/jW32qjphQGIv7
qPIGDe2IjJFG1a60lbpajergQucTzQHUlBcy7WXjJI3l4zQL9NvSGTGZPei8LCx1
OltpxL9Rpq7dBcgEe1beOKm5V/1HkxJo2XbGVcOn00GltaZkzeNYEmwMsnNCA+Cf
KGchRy9IZC4EdsDxZxdjCnRZabGpBj0jc358CVi3UlATzuVxKpYaqw8zWv1HTISz
N4ZGm4zYRsM/5tzwgN6W7ElzWlrTcHUaEwofIyr/7whkBLcVJjKDdzh9F1coZvOD
IWbSSr7Y/XAKpv2S6nSufkr9gEAZQEXE0BlD4/WTF5f0f9keVMOYP7f7EN4UAUIH
4wugw6KHP+Vky3w3tXcYdEhLD++5O70WC6RJWZx7xXUhFilOq1BFsz7Ea2ZuB8XS
17fs4ZQr4SGlxLLtyL4vD1wyXJz4C7D3wOb8iaWoEkJftbbKq1fbrV5P4tuuMsNd
iONMTOgufP5blzLKtbinwy05S3Ll5DN+YtTg6uSLMS3vgEHLUt0N5uARTBMzFl/e
//xEmPaI4fXgKlJY/GNB6y1YKchqDSsBoLuTjUX7h75caQo05v4jLlFi7iMK8Tf3
H48zej7CIw1vSI5xwU3AS3UeBOPdhG/QgeJb+ykGXlK1BLI8o7zdKEsnM8bogBww
7JB+z/Wka31h5UiUm8iWcBIDBicQcaFBTZENB1/gX3Y5jihb7VdFYW8ri7iVZQaz
YFmGV4pZ4Z/Dgesx2wXY429linTX2R3b8ciCEowTUdiSwS4ujzp+mhpuNvYkJj6E
0Rkn1I9WNxwTgL3RHyTp9Ta2ivZ9bxPf8TlkLdEGNgzsYHyBjsoycAp6qKpfD30Q
SvlxvcepjDJP+6bXsrmmxh40SO28iLA8zmqE7friS+6+4Ws5rtZTgp/UQODxRExj
IkmLtCX1cqqPEV7tcEX2LSyblaBnQjONpOEIPBLsCaAYXC0xmKDsqOYU6jRQBp09
KFFMjPEY7s6FCOL2wvf4Cq+GcNwhgRkHNFQ3ly4hXXCtRXyAaJ3Cr0Z6mgOwgGNU
Yq7W67k/Em/Or5wYT5AQiKN15+8t9igfzj4Y96bmgDF9tZ1hL6MmyOcl5IYI54/u
ZyDDcBRk+ozGxNSe6BWioCUPDdp2J2bQE2Pnl/xQsm18B9HVvRZjzx93liOPZ0JE
l9/SEQ+3gf8rBB+GWwr3N5I4207tDtbJEkXZ65HjAGMVZhNQY6YLpv7WVX08huCa
7SJpL4QDUIIb51yikhdBps061Hr4UfQGzfczXGoaqjSHDQbqYCMHfQy2HTpF8qfU
/lAx1poPjs4vFxH8tyG4hLPFckPegdHsHK+u4eSA1ECQMP14X0B1c+AV9i0JZaR2
RvmxUa+pWF1FI5JsHwoNjUQuoO3/GeNapL7wa65ZIgphEE7nV7DGYucU6CtV6VsO
0jpaAs91bYyVPCUOJ5dc1TVkJ4oNtw2qc2CIsotQjSIKBE5D+znbv2xhSEDWKHhS
wSOp5Yh3gR9W+sqzJFe3h4l5bh4mVyGtalyk7JfOpTA1U1JmTaLTnycWhAJ39kn0
E2d9W70cJ6g1n4cQTw5GMu5xohg3oLnwzwlf22Jm3skJ/Fe87oJ1SBhnaeus5/ha
PWnkVuFAJ2pdyRx58WUSAeE/lNAtAnEdjMkLLXWSkx/EZvgqM2lVWlvdKMgoWyZZ
VEnbEmS0nhIUZsieFL2DwhQoLWhs9urT2NS6UPIj4PfmFzXhBiWY5OtWn0/vKt1S
FlBwNRzomyefcNbdCA8zIBZM2Beu7KMOfXWEKkrUOZyWNkTWYEeBFBpQceraQ39z
Go+LzcdYXBBzSQAOh/iF4J8OXDwvPlf0zM6v44Ig6td+WVUf4bKuDqeXmrzWMpta
fEB8h7NLbb9pD01oXcFth+2kEVmaRIZ+/pIB61X+t6XhLm9O7jGYnAmO2J4YHCMf
hnVortaKk55OkcLogAoUxuSeh4Z/o9y3BjPkzqO5MghuE1fNEGtAWdo10qZM+mZa
xUXtSQV+3Ss7abMaIsZ1PgwKD1I9Pv0PfPfYbsQ3isPTZfbflfjHgeUw31X5hWDu
h84WksLXu7sjnm+oxKpd3V1KSYTAkVG5NjKu6QYCejwKeUNZ/M9QaHk7K3AaLtcZ
PCv9ocnLtRJHyzvK3raatcYoZMetE/gRlWShZXs5mbCH5DeObPKXTI/JfiY00OCI
yejoMXX7ItdCGiMFGdXM3rNSxvjiPZ0A5DVYm2cS8tD5lgcUq2DgagUil24wvRo/
8UEF0mg6w4BcgAGrm9bmJ+/aeE4rjv7oNz4gKJ7yAUQmCIGJI5BNYTUeaepipGCU
q4Ovvv7nYhRExv6cFiJUsK5XGYE6cf2LZBp+hlftDOaOXCAYEEj6tXXUZw4M8bsz
hx0eUI8e3Bh/fG3CLWA+VrVQMzVJVE7uraOROKcypT13CbnFlmAj+sQ5FV7fhdlG
UBkdgkaCoETgrXtxTHje8ZbtaOCCy9sEik3nv6yqasoyxHbxDAHYgAO0mQbtDull
14WRK9RNHmWSBpOeGWCPLzbqsnNDDNMG+N4KIsaR3vC+PCUzY17/U6WTzrwMLcmV
Pv1melc+N2tug8M9EqsFDTRu4fE+Mila460YiPCEiLzgGc0Nj05vPGHPHufWzHgJ
xprr15Rd0NyU2BdKh2wftG0Ey+IdYDfZDNQVjqrgR0s+ccNBV+bN7t0bgg7iBeZE
+ZPmJ6k+S+ITjAPdw2jAFZfHaYgH5u1pwOadWlcPqycJPn8OPhfGzcF2qPSO4QA8
iIFAvyw4pd4KR8t65HkEjfJ6T4S5cYQEUflVaGd8WpYvNCmG5xRux0+ubSliD0Gj
HHmn8Dk2q2ilLAtmQj4WWMuJaMZ6TVmlk4/gqFriBofqWDvh7mAQ18o1dh0Qs10C
GRjqIMWSw3NZ/v7eAnCJ+5HpRKIuiyt+ZYvhFBC3sZFLv94ozd/0/mdlXjz/e0nr
FlJdl2NL7lVtya+D+TFWOYA60W9s5TjlSj38cRnKsFI3ypJdLEHlFZapwYcT7ZYb
q0WhjwqyV0z1KIRuaTCRX3DvMnte8m6MUGS1pVhjde9JUPQfnA4BMbespQQz+gID
1doSF3ag4OwDUsprMw2YUTZriJKif0CLag/H5HNlif3F2zD2Xsnk6kX5oCnSW3lo
mwMRxnE32JvGkpjxTtDyOZZTVDPSwuhEfQtRFZcCWWRTcZ82XXhNqtA4sNCV0MHO
ZPbMDc51IRJYHsYPD79Cmri+dvjg6oPFVOSkK5ivGUvcM08K3Zj6wZDsq8wpY0K7
3K3bxmQ7xwAczmlKSZRLvyv+juZ8VnTpT0+1RcmiBnNAUpMuQ69HY3wTQV9UycI0
GgBluawmEIQFr1jxsY1c8a75vZv6P1Ql12pNnC2uq8zMkAUmZ8cvi/MmniyhbSHR
Cp/JVltnV2loTea4bjE2pv5s6vuWGsNmkwYbPRtJsB6FvWzhlGXi51zSuuEM7u1O
sw5nY1eQyYEdwqkXUzuKfDlwLuE4Og16nH1mlJkpFHCYHejZEV9ZOj96+yXd9wID
d5TIyZnkbkJ8X0/zEfhdQscRPcm0PHEJ93yeD6E/aJkt9l8JPJjT9nGXR0DsHSkZ
NE5GQUCntVAYSbNjJoAlWLDBrdDNk+j2ILnaULVLGuci9iooEP+XkgN0crlwl4qu
R7huj9VZE2HFbYn3C/d1XDL0Ee3W7GdCMjNInAyerF84JP3XDCXfLXDjC4al1FN2
SvoLkXvg37YwIlsRf4QAP08kDeDW7x2pf0IMAAwXvmdQ5aip1na+Gaz7A9D90vXa
7TClMWdEliTntbnPoY0xQfbait/psFvEAQ8i4bXh4vwhHOiFQiTtDSBoDRlB47D4
MVG882L3lD4ROfmB+S/wB/g76vwHDCkfzmDOmuHr+81hKhcDgLUhsW1wSTsfEhgN
lJAEJx+i2ge+pZStfju0qwiE8hQXmkCcNI2FpYDQTkFE71HyIdLeRIpRH02ZMKj/
sBsZ2hSOaBMl59vFknK16/+L5cu38JBCl0hwH9d+bBmqP2UNmWRvsrP8Jmw3id1m
DGlfMPJGqd5bL7S2sCgADWL9dbmWTRbOwBwOdrgGULErm8kqFgkA6UlBTWqo0Okp
ppIFTZPqBtZEidlT2n64JymV3qs21WTVWgXfxQEQM/5Vh0OaE6Il1QrS5qGYxJ8O
dU2YHS/dGSebbWzFC7JhmSZyUgmJNxI1umW+bxzr8v3McKzBK2Y30xsh9TKfHLPT
L/wk2lCdlvPq9qZpsLtMyzvrhDfvOg7bAdkrCSAGazFyMoYyy3ltVuWioJZihgQG
W9cZjvuPUcrRkzLqK9r74gSP7h2u2Q3gj+g1J4m81h/AyNb4YTAIkIe9r5+vWNU7
r5s/WwglW7NBX3o1C/6mIxu9V4Q/EUX/bm0hjHXC6Uwi7RuqaIGyw1v4OVRf41kY
Ut1BI8BfG7qnkadV0GjK7uVbK/Y3WqF1CHsNKBooyY8gkajqAf1ceITRcN66VfxK
QB8SG69eB1qe635hEuvX9Fv/6SYvmyL+P6UAOrvwUCvm5DSzkkakd5RDXgMvXwBr
mQOEcvkbNMwQzqZhMUWtKPkMsDJhuU8IiOkEQMXdQ1egu+vuMs2G6/8JQ2s4CVd4
CZ9iOOZZM6CLPdXSlK3RUniL/G8NK0Y+xg3OiIsmJA1tqs2C/fh+m3xnJND1DUSg
cvINBy9seqzNRQ1Wez9VId0esJjrK6IVxs398kCbDb4oLwypweJu/kQOw0k17T7x
7A+VgWXPI0BPSUGbGImoO9ty7afTypQPGTsXc7707j+NT7QuElY4MYQfkpv95ADe
Y6pElxBIW4dtw7xlB+8+JzbthE99GqAqIctTMlHKFvgPO8+B0TW7SRDHdGNlAce+
Xgxiyut9kxbUqBmxsPkkMfHRTOIqmvSJGFKFCfG4bLvGecjPfJHntNrAheLn1hqh
chVzLwI0uIuoiPCrLLBLv/DqASrVJbrmDpjSdZW4Prz3Ru35yNzAsCeROdAuFHMf
d41u/KO+5RdKGW7WlnuRkfEN+047RpsMql8Sfg5M1OWeNPgFLygLFQ5s6joZ2Mrr
FpmA+oDU3tUy+OOCC5kaJw/yCTayDpu2OEPbD/iJuEdy4U3LCSTXSjjdOYr9s1ua
WVPeJcsOt5HPRUjEdTSlPq8ubM8TEIv7lvvwbnAgHgz6B1YvgYTe/byEAwCqw3Z7
Wagadrvb4eBbLiFEsyAKqaYnt4GQkO7W8WKWM5RPSpRMDJmbpljcm/mXOSb/Nirl
YMPtXEzxiLgckdwuCUpA8p+M26gxbHETCc9urUKP2gaJX7tdKLT6bGorsQnOTWth
NN/eIPDn/bdrBZ5VRdSrB49g0KV6nBRqCPehWZwQDLe75bnXBXBX0doBEqDNhDBs
7CwBL6edswnDjGQTdpr8qQYDerN4TnYbYFGWQfYlXOqT81cpytuSI0+LI/vUuhLL
94VyufxM6+YdpLYghj8YKXyiIN8zULwyU1nWYja1kTY/TISg9CpXkXLK0rkgi85H
cqHsTbEF/skT64NgwTmE6+brmcy2a7J2l97perATbKhCyiekqzmw7AslF+DVrclz
wcet/9BoGbV8me8OyjG0iBK32rlDplv0AfNtpLYTc6oP6THjCfWPSq/usEeX/9c1
ZhA4/QJ4iFt63pGYi1wdpXC8y9D19/n3nBQniWCDaGp/Tc5ytBerGwg8ynzPWTQz
qdFjgNtXngriHaURbBKjtPo11OjAd7CQFGBFO/3POGVTsFXvb3f5GMeduX60MDtU
5zJg/sZaO2ds/Hm4/vx6Ppq2Y7BOAe1m8v7/iPbSrZd0P0OuaqYjrHUDL5k2Q2wI
dXzEixXAitsxSEaCf0Y+nani0z7O/9UEvSSasm474LuVHFvf7aD4QAB5ih6BKBPw
qojTSVSbB2R3nPhxGkm9yNSS+qmm5uKI/3LW3afcjNnaMt56Yby0Pu6+k2KomPCS
TwqzPRB6kTD9RJ5R2NWhxz6maRDRESi6zweecrLnIBwSjinJj3IW5ez3Pk9Zamto
wDJesnLJvn8w5yxtSTfXj4V93I+cSmeawsmqKzAnpdQl8CtbCi8MmHDmzsY45Grq
gsvtRYs8dj1wL6+9x0KP13iCjgcgtlioG36GdUpvIjJKJ5+x6J4J6eAx+QIoNjdo
LfE2yiCDpG/02AlLFdd8w46+eN9a4bhX+8Og8ImSPj6dZN0EeQ72tT9zUiMV9UGF
BP803SfV7JT6mm4K8lcDQfdXoOHzo0RQhj+wxNfAUecg5CJeOXJeoGTikGtVTGnE
Wd0AlUyX+Kt7AtOAQYRiob1wEnC3KgeHmFA5HLESoAQrf5uF/694LmCaxnQihz1Z
66LjkbIjVfQhRN2uQWCf32ZrW1S3DucEjteNH7oJ6PVzNkE9xMYAsTEs/z4ivuqx
1cmAP2oB5U6d7YBn3KDSn/MiFOJXYh7BjS6UtkNmtSu9xiZKLXUYwRHaheEihUUl
xjHCsM9Zp2jB0Y2hFnYKdLfALFkLjZe1oljUCS1l9syJcm3XWjWLyTM7NYLpXA3+
qlgvn4/OCfqHorytWQ/5tzlqbqGmvlP9BWF7wPT1Qdr4xytTmziZnvdSdUNrr+fM
JWSPAUbPmicEHtrrb0ckjexPmqD3jhAyUsT+FpwUQ1u9H488PRvgNIvXmPOwOI6n
SkHkK35cYIiuq9G8e34GoZSWe6OpP2hzT8VaSG6D50Zkikf7toZ2mswiqK5nHMfr
t2Gq9M3dZt7lm9pLpFhD6sWEr49iv7TDbZg9A8iAcjykeSh4TdZD078hmNDCVde1
`pragma protect end_protected

`endif // `ifndef _VF_XACT_SV_


