//----------------------------------------------------------------------
/**
 * @file vsl_msbe_typed.sv
 * @brief Defines VSL Memory Scoreboard entry typed class.
 *
 * This file contains the following VSL memory scoreboard entry related
 * classes.
 * - VSL memory scoreboard entry typed class
 */
/*
 * Copyright (C) 2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_MSBE_TYPED_SV_
`define _VSL_MSBE_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
crcfwTFUXEQ5QsQlYyWJKCpNxFbZZdUMSwbMbPzRi7Pq3GoYOTMgcThAl50F03hR
SYpLF4XF3c39bXGusfypM6ptaHH0KRMXy/OchGt2WqjmzWpVljOe5z7xJchg05Cm
A62dNtiUY2q+1Ib8NawZD1Sl12dnaMi9089ZDsuRf2odVDFKau8VlOpNK1KzaqgZ
0EzWAcdwgGw4UH0XFNP+7tl9VaZaAg6Yb+kVmkQEJCJkg+4/2phwOkHf8Mh/YvIj
i2imyFCTkly3RuFndvqur6o1nulTlXObMwwlSYPknFu+g9eX5vq/66ciVHE7cVaq
UeR3bCzzVpvOBugPxd+rhA==
`pragma protect data_block
QV2DtcnEJyk3a579yTgg1ZjdWzhEcmHq+sA8vWChazjSsUD98k0Pl2Mk8Xnpf92t
gZUuUUf0XL0Omt+eD/MFbicBMd2G/4gLW3f9Hi90QofhjdXsuHK3LqMO9o9Jna+5
L2lBhUqoee+5aD1LVsiMAoliDf2U94w3wJncD7D1SHOjfSe5mnIhnTw+TLWbayuB
dxX11SXKeaEaZ8KQ8d0bBME/d8nQN78G0Z5ItH2CWIXb6X5qsd1ON1sDpXrv2r+Q
WglPhfE68rLFQbNLvPjGKwxzGwSgcxOZdcooH5gwCaA17mhddeASnT/klerDtC9t
8f8yAY2C1dmp+KXd6pG8XCplNCy7A1H3thCntpBPQF62puH5iZmQc+YRh68LelN+
I3CDw+fDiTL9n8ujASOVhInNg7eCQMmxEele2EsUfQfw68aLWnW0XXUzl6Y1DYCv
GIwPye1lSS1DDuzS2k9l3maidx8HRpG6tBbHXkbwjCuWZ9ZHO9DvfsGNVkEbRAnY
T8z8r4rHb6ZbXYrH2I6EUYZ/2uMvCmaKY31bnwMucn6vWpvJlQOZebvhX4FgpIIo
QjyVt3AHAaW0OVM61okjgNe070yRZYIksr58vhZu6iA7kY21GKRP+cLlPUKBTAed
1xwrGlPS6aqgRBQOzxiNdnkTMiyazmJUOVA1fBa1gKzr1nGCVvfYBEtesZFPCelh
5kBDF3XgzL8x5GmzJo9cNju7ZP80eFxISdQiIF0T/3m+gb5u+cAkStePhdURDV8h
yiOozuK8aRm4cUQoqihMKCKXUoKebiJkf3Swqc3QbyhLHABj1mijAub0L/CnBed5
PzHG1A8SfZaGGGbiqpVMNGNEt8NLPMkQspiUBHJJ48ld9VLvXF1iFgxtEPmHWCVc
BM7EKbLHy6GEzFGbGH4lB9emHp+nHZnh1R/1GU1DDDttM5YX9Vl2enYcx8TxxE6Y
NkbueN/wciA1k+dDt2dy7BTqEESaFL204FM5ftMmSgU8fd64yJ3oQCpjQGIWKQqO
40adktqlAsFiko+osAis/Sk0iajpn3IYw5GAofCWgDpPT8lsb8azv0EnhIALWtfE
3X9W8k5FWq2a5p/N643RSzltBqviriKvEZ75aBsMCZylB1GopWkaqDAaCmkFFAu6
XLt6FSfWz/Fn+U3uvlbUKR6sD0tqeRKdhVhch43yvOjnyLdQEur7WWgZjkMQWYTv
KzzC9pw0bD66Fid71F6YnUs0qV7OB/sAWLekqsW950BIfq7JrVPeVRnt/vLFWQkm
5wdodmC8zT7mbO8EwePATPJoTPftntkly+/qfsd7xyRspLelGRIT6512RrLzHBNJ
OYycJs3MIvf4iMy9k4SwqZCUuVGn36QH60NXq2Ndb5lIp1M72ZTBqb14B0WOHC35
8VmiDatHoLksbXNa9QGkxP0UcLhJGErPHk6ZTNcHomwOsc0FROwWmlVArz4eRgAd
AWMgPDda9618XNlTe0/IKStG7nH4IGQU/aRFTkPVs3TShv+k1oy5Jd/hElMoNNAY
KySMmBpodjOk52ZctV66iQJKRyVbzYPxTOmOl/hDruNy6JwM9+VqdulSeykorJ+5
aH/4BgWlxan5ydWJBW6HNErZ14GtyTl+QQkUpJaZUTifOhiHxPuQsC7glYQl45P2
0+VVihr4Vox+GqL9i603buV8/LE71hDZDrFMOTJahYD/6ApiHUi6q4EVQPGNhquE
Q91pz9HHypR+aHELbu1Fk+GDfjm26xTwD5AQZKJuBFY3kW9bjDEng8vUCPTaRYuj
4H8VffhMLkTBN+nMDC0nRlhnXfQej48jdTYPw8c8Cnsv8LKMp1IZ5Uc78I0hKM3A
yver/m1Lv0jXJDDuDHqf+NCfiWIVW3IwZCiFNLhLcS0HjnaE5tEyhC7yRgLclG48
0c4VGW5WfwCv2O3JNsDqp1f077m6e5CvaR31Re+IUwfAdROc+WqYi9hTCnXYgOr/
OYEvMv94+3cDaEAD6UeksRTpwTHCgiUsceN2VtTmsJvQ+YcYYgbQXnlGKi8iW5bZ
Rx3vFMBn8jgrGQRm1KES47ddHYA7/JiDs5o6YXS5HSFl6nAfvzduDO7mYGrIVg08
g98IdGJkMXYV+lSx9egxGvtjjrnea2TenyEII9mcpyfyhra8Q2Dw0Io39imdkVRa
wba7jkDZFFOYW5dLDADpcZYxHmYUgQKmwSbhCg2Panedar6sHLg8ysi5bbNVs952
UlZ1egjR9jt6l6+aIYg50LxXt61sijobHJrFr/PsMPDEgUcJ4Qpp+B4r4485izdL
U/1+A2W38k4BNgUtwdck+hfZ0eteZ72+CiVYNYjzhzgAKV5nedyMdT+2BcW9z0Y4
U38n10ej6FadEA0kmHGmUf8G7LpckQxxU2SJ7YejCuJrV7hZ5XJW47qmDEG3x2Fk
qgGxLrgZ43Ib9CP/9G2WdEiVpKkHkVAg/uK671poKdO1rh6fRJ+s2bGuXD6EJjpO
QI5OP89Vj2bMHFzKc/V2g+aIOerCIba7/+Luysa2V1wgXHJc13Li4UR5hsHkBKFo
cMbJ3MDN1i0OvCbP9MvRyrw41pg/wxWkKD/QigbqnpWumfaGcKb+/HqJDS+z2cMb
02X6hV+UuYWM7+LRdcWUBpHMWcodJvq3L7cUPzEABlma9BkSSQYgx5PWuVM/nv9t
cpJuB79GkZCa14ZeQZUQa2XQ9UQEA8I3l4DOTkfrOxX2T/E32LlA0w9oiHTRhAiY
cyAQlkO5MAkTmlJ9u0uqoFqXw1Ma4gyLBNfwGNhPWjmOFYWDXQ9oX/QJNCj3gory
lk21+BZZnWpVk1HtCw+hmhY3F+QrfJb05WWX26Af+8g9KC/fdZQy9+m4s5SjqKU1
KSXx8RpBudqA2Mq1PM7Hwo6rlJbHfLqUJd7syFoL9bxap3K2TQHK1osVUiDvswDy
t1TGzPU6stz4el0MTEILSEiXMQGdfqVaUyGDK120G/0U5EoNsWf7YurDNVEOFrWD
FkZdUK9nZnFUivKqe7Nsw5vGZUkgK5A79Y8Db4s5rPEwlksdGSsZ1JF/iBQiGf1i
rFkges/ZYSTp18kllozpYJH/mDZcSZbaJOycePGG37AuLM41Gw+YyP4L/pulDlyb
ke5SKkUCbiOn4q09fBxxZdOM+CA9lRDBLxJ4C+WYjk1TqmwIu2/WxMMM3h1VU3Nc
gRSgAfSS7oKy5hXG+Cg776A/IvEpn4hZJEA5n9ReUC8RIXIpRhAQW7eZagLYxqzY
oOjCcFvazTlel9V71qmw4x9aylicluraaxTdLNSLS6DBefQMJFo6w8ja+TeA3GOv
laNNG6mB887aRfxUIIt5GlPJPJzqSf5AiNPZ7W/1eBxeKK3lLvhE+BFK8HAoDuWC
aq0ySOpu44zZ1fCFTjmL96RqRpAubHG8Zb2XInwkIZAWXJ+xSJkQEVGK+4Fr+QZt
2BLJFZG0C5hPHjXCNhY8vyjuYr/vqN0y4jPx3KWpBZd5CGgD2W9Rg3qnNTIqvLqj
eb7dOmrFNNTnrx28rTqX/1G2Tj4tgY7Q84cs5VuV6yfKtHXx0aaEt0aS9gYKeZ54
oS6u7+CsGsutPMwnWTYQxJMEQRchxCkayFKpUZ7n74KGsoFK+pVNSL9+9NboX1E2
VODf4M90QPdaNg1pJ0rKtAsC9kJ/TgqDI/ABi/tf4Qs32yomZyCoVgdPb8rKNpdF
u+GfkzOopHmjUDnwYkx9cnXip1bROPwl8SpApZ/eBs89B6mW59mWT+k52eiuPm7X
qbSgTFNZd6G34iBuZsouajYgYTsqXT49np5yERZp3B/a7PhqZmRrWfF2xFZX/OrJ
hexeI1m9yPRubBSKBOhoOt29cecPBEx0ee77jQopjEDqFqng2TDqJF+CXwRxD2Lk
oQbyXqAsE3L84J0FSxst8u1DqYXL3PMA3T/agPCCafHEk92subSnt4fCww6c4AgV
vQFtvUneHr1BJyczeT1n13WNOjzD2ljHIl5VWftj1v4LR1C/6qX+0R7SXXJ3uG3S
2qE6UXP+6PP14c68Q0a0SskJB2gnPlhuECc/egn5syHlfZuEVF94+ovL4VbRc9Gj
3xdA3FeRnQNvnMIzif7ggBnkVMPd8XUNDE5tBhd/sqDEg/fO3yLMsElNYof+mExA
m628I7Iilp00VlYcobJfXSVnW+v7IunzY0E5YpoYRTnyNiAweUDp2GUZgXHPrwBN
L56I/GsOLmXnRJWqw9gfNaeHhdygRVKFGA4iZ7SxZWYA0ZfcvaIw6p5MOxi8EG/f
8fTaEt8ECyo/Jza9axYBxoVxLRuqBspEfJobxKuiiFKOEG9Z5etFTjGHSzVijXHI
/69pb64k84KOMNaJXi+u7hSk9BFx6W4n9dvTQGcQiZYX85/uBefjH2me1Xfmmqye
U/sesH8h/4kK3x/0JTQpkTuBCk0d7Q4cUizUSuAqRnOdJu79VoImumRjnoTmKv6f
0igCz94KbR5DguVj3Sgn0/u3i0IxTJiPR1SBlf5HvZVSweJyFZuZ7+cbFbZTCNGS
PGDNS1A4t79LaYtns1H9NnwyeOTkVh95WgfYWTS9PI8Zd+AKBdxsSoLMOHN+KnFi
Ay6FBCfRU+nuw5wLuR+vuwli1EbqS7OYIxAKmBZm1CfqtPckoUpg+F/mJGwr+2kE
i9BWmUocMKS1uwQvv4YAgLOgb+cUhgVW3pkpMS0bxop+wSSDm16PmPCidW4k6Jp7
ov7f5FN+yNSpea5HRuCVQYmQ/lmttR6dduDzEKTNu/uAd/LxutyHW+2+wZo45SoL
Y9en/Y5DA5isJNgjWvkqlBOruGYO1FRoDBvK+Ay0Xtl19Ia5ZsJcQ3LW3f7NfPjC
ZNgs7vAm+hcDeixaNJB5qAu4g/vUofgT9EwoENoov9QOsjrOJqsb3wVo4oCxXxqO
BVlXM30R/T9FjWU73qWSJT7wePq5xFja8nVhKAtQ/72AtT3gFIpbZceStn/A49zA
1IkSpIIzZiyD1/I6ATID584wWXe1v+uR8RM4WvPXElyLzd6XZRgOY0ofAXl2ix1U
5RSB9NwWHM655EvaNhUf/9xxPbx2EkC01HnJgdTAlvvG4KiXbko2ySuTbMdJf28r
aqC/KMaLBAEVCQb+WnKB7Eromgyqm2U+PCOlZdSwyVrXZCd+vDlcI4IeeBkaNxPj
o05afggrxosRNxhmAJCnVJgGpTJtUph1UHNWhQSJvLRjTaB/H+8NvmZM2Kv+SpUh
atbtf8TEDIYQG6EUxt4VCzUAHo/3ygu9tnFp0C+XCeGbQiee8K9904IuJW22xjdN
QMxQoCWMGBbmgZ2POeKmGsmnYzDTWdaewHHK5vO8eTqTybPTu5rEvTVv3TnQ3/L1
m0vPdn5rrlaztsTDEwFPP0cm5R7HlXAKBpDfT0rInMW6N2utgNMZq2xefvGUXt+5
tguqo+ZiwZrX9ZjHzkuM7j6zzsb7rLGRq4lGaIZQeUIa1T/uyEKZ+A9pTU6OA9Um
inaHl0hqyJGNMBszlkB3eIiZ82bXBR9gzZvGKZIjiyumslDs0L+ApA7PKtC2rRam
oYgVvGm4Y7v6WD+/o3VQjeBnViDnvOZP+vC72HNLQkY/ST+8rrejtDTMm9qw3vI1
4192Utk8WiX3fWHRDsr6DyTt0+0y2iZu/QMHkUnBtd0khbpTPHzjBpvIfMuPwiDD
Zlwgix9ObVB6iYdRjLsp8Iiu0JRybK+p6t93TDE3uYgwTZ/EKtgaVeutq4UlzWTH
JgBW2amYv2W2inwFxqskRyWgaUqLxTXjDMBtWvDK+5gihpw87+hPedXgVlAoYPZs
22RbQAG3Xar7IQNkNFB/Tz2aKG2Qx/Ed3jjbxFR1CtRNX0fSWaJUVJpq8qRPsLrU
XJm5+X2g2AdCV6WWB+G3DxsL6CmFvnVHQQe4aw4pUzbSlgo8rGvFJsAjifTN0lnF
NniW+EEdGta4MS0HAstpmZwVEMmlYoTF2l3r6D5IUKZM/BtZdRxjW+XPTr2SVqFo
Y/Q4PiPNLjI6DBNqsV98co3e5rseN8O3FjZOLAG9D+NpNp62OlWnt9OesphVKIUs
xyK+YiLvh4PUiTKXKMeoZx/qXlCDIvYd8Kxb0Bt7YHwO3A2RPVvIbHyF9V7sUYa6
0wQz3OHyC0kTC2lTJizDrVBw6viq8h3m+vyuSW3G6OMPa9hxP0ACF83O/5fCjWb7
4t8fPDgkjzVK22X6vT8Jtd9UURdGUjVzvtPrQLUZkjzMH3JwqW2rw0yVcyPY3NDP
fUtIpqNwHUX2lvz8Fskaj3BLztIf6ToAbp1uVewquFxK2xMuieHycnJl2DiYyyh6
1SjIdfo/Ul2PR2XM5U7WB9tJsON/gqhVGG3acFryRWtCceAnmKiKpX6RLZ48+f1a
/NCbzorD+Op5BaIHQqCnurfb74Hp1FTC/5yzsqCsf6gc9qfg4owJRn5mZr3XIP0N
TMYYWJp7GA2DvZ0WBrfxLxjhjrwJUGi5WCCd97/cRs92YOkd2Bb4tZLC29238d0T
3mucjSOH4jToBKwEnUqsNaeYbUMiC7luZ58VmQBitghlNRuOJpvMDiyqcw6wolQK
pxXn3/rPP1kP9IyVpPgNqzfjst7zNkydrWfq46w8XOC6lGifKvns3q4f3E0Z2uN4
5tkLQDVr/jT6+kcBq2SwNXmlCYBk/2pNqqCxiK6LBve3bIxr20goUMSkWzxRf4lV
uyigSwUnJ46u0BjMytjby8xheLnK4pduypFx90ao0NWr+5dtzoQ+lQV3fN5KCWlQ
sSUAlafMofeBVjkqhzranOWpvAOpQzKkpkKojeXfdxWUy4vz43TiNn0hTXO/3qzq
aSHw8GmeLyV1tjkyu4YXhxI09AkLzREtwlNpfOd7Q+nQoT9b1S2fvbK0jlZyYOJe
5K7ZgtCEhnhKk7pIhXxorG8o9iDQfzaswaUssX3393anT40GRf371gAXPk73H2dt
OyY6Z1gnrxRruQnDB/j5A/Q/QT8CLDs0Ut1w2oQJzGNwSnf8WK2dbKd6DkbH+Wuc
AFNiE3nDdKcdWKWDtGAtFwmhEQUpL6T9g/lDM6JHjK9QlWLzBdOhyRbsGL6RKdeA
NlOdMJFC8gkSbnfnFoVgTrSVdyI12/T6b8kIylv9aNWQhclqmmIROuOd3J2xfP4k
PZm/BgFKn4VTnIGCa1MwoiV0jIHidf804ja13hEzRZvv76VCHfer4fHI6igdf1R6
5re5LyHJfUO4BfrurkhOc0k2kCNAViwW8tHSWRmq/WjLtePxeGzb8eGcIn6u32mz
OcgRmKCI90YivON92zFUEAtOB3HuQUic83nNEj5CoywCnQSAJm9BeOWFC/Qs1tiT
xvuKUJwlikzimW0mp2Z+2BRsC932iZPUnVRhOGyAyErQCzgC/YI6p3u4TOCCCc4K
Kqxw/jBGgU3sAWb5eaghjDT6JNSXkpTPj8hBANtsn7zWknVEr3c2TQesqOTmO0PC
Ti0D2RtAorwblx+ro2pAjBMoLdU/SQXQb7Yzv2TEcEb/TP6M7U/Sc2CKxkq/kLAY
+5WDyNGFpYMTneCkENXiVZxiSP/9UIeXQjIZ12VA/mn7Sc6OjxvO9hEdGfNsTDjr
4HXvoHQrgqXN2SXvD0C3SHAiPKTNGiRPnIzuWJAD/XXf9qkDxixSAJsxv2rJx6wa
IFPMJFz9dE83/ZZN+ucFZjYe2Itfv+Q/zuU9wIdSIzekoB4oBSRNG5FpC14UyFNr
vtNnVOkXJwn3uMkly9SNZiIeurDolDffazy7fX7izJ313O25eiJhqB7pfjeksoEQ
vOP9nXu6cwhGT+mWMYZKE8kv1cPKothqRWwa0nkH9GL6QA/hD4l5mZQAUn8/LZhC
E3jDQYNNJyvdVf1d0P6M3ae70CZyH2olwareOU1bQlAVX/dtvHwYmnabcnWi9U4K
RoKflEkUHz6sG+XFLWOm/Lm+F2fYjRWjiZWQMaLULvAL8qh1zF2RO5vUNfdrjmCw
g/cDf6eXQXgwEeWKkwesYq7Hydjpfuj3KIDcVrA92UpurRs+nOODFtD0hmf9BRHa
cKlApTLzyaf94iPHccetMWpF8yrYYO5q4rnF/CI7vmpGmoZdMHBfKFzvD5e3bVf4
CuMNw2zIAAcn1WRuVM5xwc52LCBKHdqBcszG/w44yxgxMdwYw+S0Q1dxL8+NFucI
vTqCCW1OOXJcqKgrmvmZttAHu5ZX3CnzH6kwSkWjMdC83xlTCq8zsJPoRKHo16QK
hH6YCM4WdObE5lEKS/0o2u0+o4BxIaFwXBIXq2uSXGiyq+hi6l17qXZ5UGG+yRpF
S5saDEKKkyQFEjCShdkU0uXlp2ct29BF6O6Fgn8ouwZTPfuQfgTowQyYAv7a/Gwj
WaFvmxBqF+wAS99mW21765zJ/noDO2Mf0GvkUU/AwyxqZLzyOXnRuTKFmc43MOjq
CslSfb/ePZVTzBNsgzyfDgR/rWN34/DlPZoT7oHHd2DUj7rBZondI7FPsHuAaSg2
3EY31e9GvcTdvxir2yH5Vv1nbXgCMIubSiHNwADFxDH9RckXkM2rgG47dSWzTp/W
CFW5517IvnuV2hgBtt9y9RXuZTqCf4TIGnHJmz1AcuBZw+0YRjNkw5p/zoY+nkRy
Fl7v/ddvCDB0+2gGghK6RtWhNKIm+luCCjf//4SmIaoweJJpSdfqJcLoN92TdSug
i6zhYmCat4XNyUufZRee/t3KmlDhmLBUVE4nwdu/G9xwVyQ6q8rruLPb8cEMTNAd
NnBIehoTmv5uOUDVJ1EH7BTo/K1BRn6X98yPXD2Xkr/Ye+WbhCphkYN8gOflkdXh
77TSk89AbMVnw9itdgejm4ETtsBmW5mLOQICS4uodQZy8buvKzIipF+D19mlWQST
sjPzcX/6We4rKvgQqew626XRHRcBl2ZM0Yf17UTguvhC2n02Ozf8zvfXyxFnGPi7
qQwy+lw1oCJin9FFRPYsZWRGsWmz4dJST+f8eTDM/vCbmepE0f3j1LgeFHGVXFrw
pnQifZ9lH08Sqk4CAvQOMJVNLP7HVC2+Zjy2arPZnenIvRzlXqymTvqOT7l5gyP8
mLbKY7GDmoXYCht6LV1CpXHZjVzmMEbsGNJdEnD2+57xyAH2DazNx7LrhT+CVCcu
LoHW5l1btGCxBIQU7FKzBys10qrGU+NJXev2jNQP5XjRbgvpz2/EM4RGuzqU6yUW
D0/yku3mJV+3PS+ZJLhJGJb2ZuY40/xAiqNC6wqoZhwJ4+0mBoWEoXcWNkqbdp1E
9n9iUcdeCEgdjuQWIzRHct2V3J0RYRAB2DT/YNmwyhgATnmmFgtiKGvhq5Clyk+3
NMveFuG/XqY6nr8Nw5Z1qiqgDgcKA2QFp5z7u8IaEm5A82OxoI46QulIy4jwG3in
o0/tth4YeQa2/khPSVRh86uOnU2Xjl88O+ovL/L5p0Z02jDak8VWoV6zzr+bx/kM
8KyHU4bUjsO4kbGe5cfMH5OAeZRBR3nfuNJNh3rsNdmk+EPaFlcjsu6rdc7y+4Cz
hXDf1yZIQnNqtIqByGVwcoZYjzIQwTjudBWN9yrOKz6CIM3jE0lSpHgqJQUX2M3r
AX+BcIGRY3Qmg0A//hAxegVR3fH48rcR6EaeCME7ccCslyFICAvYgkGCtBZARxXV
Jtauu1aSU9M9jVRVtXXfvpt8tll/kUUH8b4vORcZfC7d1zwb0+w5rjEtIeK7Fgxh
QhmfGZANotAZSRE5sYiHB7TVvPm7elqVLGP82fjv/N8IlCTsOuQQpEbyKIFZBHSG
01O0ik4tJPIMM6wKeinWNEP62Bvrm+T2lmDCBg6Ub46f44JDlJRq5YjDfb2cw63N
0ZYnLHjp7Xd/Ds45YlsASzjyo2jmGuVsBezA2wrc2mLokyh5OjsEgmTIkLDTdyGP
ibDl+YTi28PlXUzJtPx5kvM7d0J6K+ZYOfO9AdVVIblxDSfSzMPZDw3vG5fltyhj
yypMC0hIyjZoPNBkc4E7OMwZ2XEbxOXRj9/UYp7mzt8Lhj46IcdK33D8H9awVmNw
McagZjYb3KAwNH8+3id9XeF0vHe0FJK2++i12taKzlzR6CwsQr01XtvVykCyfe+O
XilNEqm5XbL/s2QWHmrc49vLtwPqZuR6e0aSplfPrfytMV/uiJMzkqrq0z+FjWcb
ypIJXeul5eGc5uJWGHdze6bpdjE2kEDyfVUJo3IYTlwKlMrwI+sm4b87JIwV8L8m
cRcFu6BQ852aBfZ6WxjmaAkWoZoABE6hytsVpwOZvHD1yi9EA//eIf45KA6MocFN
9rWfF1p1o7qq90/tXJOionpB3GMgD0IIzJmlCNZluAIqgk4+XRV9NpEFS5fi8ihK
NOq0jetkWuAIxgafI6iWvr2m1SkjmmFSSXzu4r2uYxXQ0KqTD3Wz18Uqm4jifw9p
N+dniSt92dziJgz6a04bLIgDDV7x3Wv62gWD0WmeT79cK56NhYIL36C04vtLiJu7
Zkq4Gp0uf8BvdCPIwNDtyJOyoa4Q+70wmbqUt/xUcc+CKUXjFS9Q9rg5ddtmQ7hG
YMUC4u6C1nRmOcBArNoFiwYgpEdHCAUjk1SMOn1M4uwp5uSxBGHv3lOYr1Lc1D+O
FucUw2r/ZaYZBDAzZZRTUMznVHRubrUq9IP++CCAV50TAGn7yM5sreUau/NLtu7V
Afyyxvd7pM1JAC/COjrBDu9XyLKkY7DacRmPNnwQKh9S16n6xwniRMGrcbdDz/1G
MBB5zTjxCyKuLvgnq0D2dugzK5ZBinmS9CxZaWA4XgdwRdez+OVbHUsWNyu0vihm
YqJZ6UjrELYh4oc1G8LZrpxtwmZG47bTQ2QePJAyVr5IFlP7MtcNaVF4JoXhSmoT
GkiBl6JEZR/bMhCOlWsmuVRrT6kq+1QrWoonTFRz+Wlc71WDuOAlKia2vx/uM46i
bgh/eWXNwlzbFkDne10yWJjmnG9Wr6SFQrBSi+WGvpJ9kb6kPLPUuWhxXLf3/Ofi
//+GVOtJD4C0+Su8E4VAzNi/g2hQOOjGxxvHRVMCsTJfyPuvVYXj0sZVvvOyj8F/
GasllENrk/IVI7o6aO8jvwEnlFvR0vnRZHhQLdMfj/rIiUv46f2QcgimotnrXWD4
Sq1TCC3SXTCObNuKa/5nNFb5AIjGYYQhM5qwzZlAgVudrUdg1OQRzRsnY8YgVPze
RJMrG33bsmY93GGUg/zzayRiiYAHx92zpBzvuISdcJwqmWNnzcn8pFkOjFP8ZdTw
UQ5n/LI5exdxx8woz6JP4BvosrbXj3CChoY7BTYOkL2giNJ/807ZmefiF7HBj95E
0x7+DK4z7yuZn+e6KIfu7BX2u+LOXdcsG0RA1n1B5GSVrNekM0nuB9r/oZBG9Dry
73uTH7C6J1nbDDafyQdN3cwH9eGzWQMCRCkaiuASS/EVm+VH8nbQjZNpjNFIg8g6
cYuAXqAF6rVW9jXh1Nd5pS55NlQGTLaTVKiaPNcgNtGCN4hHpuJxZGYINR1b+e6V
/DgfttLpaSJjFnPDpnyHdJg8HXTLMBdt94RSjLWZmThvtdhCnK9r/9q+GWeFvjO/
TqHpJLjFU2rRclDptjFviGkCPuU11YC5jdOwOS645O2MT990qfrvDN16rR33lcjd
Lbjf1y68tOQimtXSvKUEXoPxRgFXX9Pk1sguyEUvMX8FiX44iyfBGW95elgSF7Bf
ERAQp6v2c9rhohOe5nBA5PAPugfS34K5hNYW5V03DeNJTZqpll9OsN3UvisNht3Z
p12/4cHOxtw9sexhWiu/iZRHBFGF2LUy9E7pHDBw0kxNQO9Wgwx0fCmiGtSiS9+3
Npedc+Rn1OGsJVNi6xmb9y36BKGLdUdG1dp/1OHSbEur5i5fMAKf8/q3W/yT3p1c
QMOjRdeUudBhuAKqw69EQX6BvCOMwedg1U0xNyepBGPp5I3RukuKHQXZ8SuihLVU
C6YZh/18AfxgKt/L1dAey850Y1YJA+Tf1yXCj88JyfVxnhoMuXJVt+BPWW/an8KP
7sGGqtCfsPkvxDqi955ftV0Z+AXcFV4M8FSeAIYlhSIqKWLCXvzjR5xsEyX5SfU8
+q5nledna+zpmOlRTRya7UfTNMrEa6LaihdqdoenTQ16F+B1bHWjqJjxFjptTbNt
l6WgzW4uI13YNccqzCcz280vgOJz7wcfTYkJNPrOFKO03CcQ3AGOftGPpiWQ8pgJ
MLPTgG0LlhGDYnvBUcFD6erxl/HOGxLD38uNIK4YnssVoyIFcWaV6mjVKBkqfZHH
cZR5ZuUZxWEmUKwe362lADLeVxpyZVXq1Z54VXC0TlNexAk3JDCjOV0arrO40CH/
Tn12sVyUw4mZ045HphC89ZoPDI0kGV1bgm6prRQP40mdklHM3X1rrQDOtxUjvJND
na/8XFE9yDz+ReKoAIEhWE6lKtOYITeoKuu2nliJaKoFWhne7tMd5HNd7l5W5TkP
GOv+6ER0R04J340fGboOxgH1QBw8r4rtsnEIYzTjffxe0z0Lq+Dna9gkfpyx1mvg
3nk9j/Jsx72PkyjXTMSl48HZsqZTYqvDiLYUkctbv6LREfGyPc3bu85fLabQ0o/x
JjccYU/firNlzc13p5gAap2DuIB/S6U289onPMXP/1MbhQ/RojqtKirgD6rGGyAm
JBbeM1PtVewV9LUBYwR7c1Tg3/MWghvjt3faruACj0+Nn7cdl8syvRS7Mqg/VHve
Vfaysr1p5PKDpDlWlkwNOj8PBJO9AoxBtrEjCkakm4q3Jrwuf1xqyaEr2O9Sm+2h
oszuMBpXfLyLkNwhBGwr+WOkp7mFxrI8cwiu0H9Va4qRBCPbbvzxU4nVlhq+amEq
UBk5BVw/md1aoWHR6Dy9AXfZarTt+czTDJlVWBZmcfSHaICAv27y57PSRwHFSFsh
a5a8mDcpuZ+LYNtXBxvNQUe76YefB2rb5lEGLggFqM71iqd5fW1X5bvq/HXIe+0z
CSnT3TJg9bJ7epVULYRNhDLoLqXNjlbvVXUgXQ/w0gNJg3phao64cFXqfVPkihzZ
nmt3sU8pPxhqZU/y4UJ3e6VEpRph/J4yOX20Dluz63gOGWUgFIjwebBER9BJ46EJ
Wtt/syPzEHpAHYqNq4JGWdkvCSHu1eVh7tekKJTOig897QDZX+GONHhgqK+U6cMY
mkzxo3DQHDFQvXYQMvOuMwWmwD7k3I6fBZp7NPWJR4WXHGBI0fp04Mt61dKeeIbC
k5uDdbo/gZ7LrCnzcQ6t/uKaXq9eLk3Jb8MJiSDKHlHWC5dNxsfO+C/GRxxIlhdf
LACNmxb7IczxcPrCaqwO7NmKzS8Z/jvLUxpGBb4leOE3JIBoqiO0OLff3ioS5tTN
2YivJMwansOjkZ6bOLujt/uz6kA4nShCqSEn1iy55xVTktr9X/OwSsStF905lkuQ
d8bop2ValL4LLy6hjh2DtKg0lus+uvHiPXhUY24W3zXsC0iVucYoh6YrrAb7F84I
Wao9Su6gwdTjwdP3sik0kJS41LWKtyRP2jsVyivkSrlxKHgFeOU/vxSSBUHEovkU
RUV+dCxrQt2Y1iinTkmDxx9fYR98MjsrOGus0FUA9Ab1X43rozrA/0lz2l4nBqlh
5L2HSBDFQS+FJVdDwVu1f3tBosf6ja//ikMJPTH7ZrNYVzn75WqPhYaHnVqmVqRK
x1/S9Q6mlnAp8eQaGxCKrDaiblUCMov6u464gv2sZV1cOuWJ9ZTu4mdiPXbA0s9a
SXkv4WCCJyILdJYiAAcxild5my3dVi/aE640NFDkMpl/f7+2Xr2R98QeBNUVsYuV
DWWavllhHna9u6p5J0GzsaodIKysNRaipZbJy5LZKqc/cECYcMhE2lmWS2gmh4Ed
U+Lcla2VdF5npdVpsF/CDesX9zTV2qh3+CF07zGCz6bUlbPMt+crDlUX2TUPpWcS
SQPFKFck/co2nzKQ562yfCa1KvDg9Bfo0KJp6+v+YfFzARUUKf3wY/4KwJVOLLDI
Z7JbZ8ToId08NlkSurss+4UHYwhWFP7EDu7jvSlX6JYJmkvRtc93m7T9VB9usU2u
jVv+udcwdWOdyLqaI1FFwAf09Lbr7cECzApFG4shbcBnbKWEk8EKFgE31hDEM0FR
xDPKEQmXWPgyc2yUcw/yG4nrq75Pb/JaNF/BoVCb6TuHfed7ovO2vjF1bVCrFHMB
5nSGp9u7EkaZhkv7RfnqSiLDAOPvWn8yrKC/s0afpweYJ1uNzUNqI4kw7NddBSGc
b+/trsUFRXffD2pD7JrI/xwHz/1FwU35bWaK8laWcbje4Lt/CmuTXFGQgOSOPZrw
`pragma protect end_protected

`endif // `ifndef _VSL_MSBE_TYPED_SV_


