//----------------------------------------------------------------------
/**
 * @file vsl_sb.sv
 * @brief Defines VSL Scoreboard class.
 *
 * This file contains the following VSL Scoreboard related classes.
 * - VSL Scoreboard class
 * - VSL Scoreboard functional coverage class
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_SB_SV_
`define _VSL_SB_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
oswLjUDAcGF4aX+0AzW1veR5tz326+2qeinK4Q8mftNhRZAmtQEICSwj9EotTWrI
wlgqQrwNgkQStknYDzg1UEPtxHk5rXAJ/58JycUV/hCl7NkBk9ONhVw/lfufTjcF
1vwCwj9m7QnD02wGwivc3DJYyRP6qei7DWiLx4G+J3oBXmZ7Cr3ts/vaSD/f0hYi
G+ilf5rsvYYzQrfMSCdWLIabjLhfJvZjKk1GpDaRInlhpf21MMrpadvGvZRxYtUw
38aPO2WYIbzyG3gMgehoLIINZGYdYDm9ckMbnm3nulienxE8gSqDx+JDcq3cBo/y
zHkO1FNANzNM5Jvl8iTeUQ==
`pragma protect data_block
W1xGKiq8uBwFouSGWOLn1TfjlZJx6PK0rrd57tlWG17YkFLXpX7WRPdPuaWPU/tR
9KNe531EUgHSOJ+kCeBL1SYJg5F94LXUYp/8/jREj6z3o5Qb3RVPMZQhUjUwsBpu
1k0Iw91Srz9XgcYLhINgTmOud/G1CU62GiZ/8Vc2wdM69MXEHGhNmhcP7xQKN9bE
YWUd/NZ3gVRO33+BQVcHJZSlXkbA5qyw+yfZgqFVZbrBovA2kHbU022hiHW2+Iva
Yd2Y2FhnJz3S2tExx9rkBuMdJp//aE2m8ZqhaNv7QT+oCu2Lh4ASjM0yq3D8LoNw
q13hGTrjyeRkYEoarhe5YeN0bHXCXWXGmGm24DMD1LWyhAsANgA5FScdERnrezTS
+fxW43mlQGTGEjFOpzVZy40BjCM/kzAPMPkRPxn6tsEjJ0L6CJCgIP2N/l/A53D+
zDT00rScbcX38GswP7QNGwx7l7uoi1y0jfDr9SBq/TOSU4NiNipaF6H9ZFWsS3fb
V/XzAYv5uRB1g3N+zc/w9X0SXLlz7ssd0HcNdPyLZ6Q7sb9tRgwOvRdIfo49AQKA
ytK6JFp2f5bpkOyhNwE/b8vzeI6v9LA+5kfteAq/geEl8fAfQRIPYkgUhVPFHS9R
LmJUjf8ehfz2HAkH3iU7V/yEip2lGajBNenhOEt/jDt3KYgjFMAN4HzRtq2htZvI
mPk73f+0Ki+17MDRqb8zjbHGgd5A3ni3NPPnFj9rE1+WMQRnh1GqF0MOGfss9l6u
WUbiDzZsSkBc2ze6umWFq1qYCgrh63yqcXgeR/jjBwRGzxJGfdEAFXFwOuQqM6cr
MYHNx8LeJmBnCB2xpa1ZkPkfOlYspklnBb/8n3DYy0J8OhIWbGGj16UEIRMdPs10
RlY9Op1FnNl4xzQmDpi4eMWrwsWgL+RCk+y2UsiIz0yvADlPkM/cgrnFdgZK1qv9
KZyA5idkh3/RDUpFcyyB0ebZSHnDdHqk2ibdKh5LHfBgCr6MfpeM4OCkPBUxP642
OeW+GXVurQR2EWSLMh4aJO1eVbJr0i++cAAwtVKd5m0OzHtXe2o9Wf8TpFqfqzX4
V1IPEFpTyuzhtdHC9fYu6xnG8ru/x9S0mGMYCI0Rm1m8uiwdK66JprOEY7yQC9gE
KVFmQFvzoMvx81NaawHw6HMBKzF+X9mBUGATfCqFaUuOWW7aAg2zZF8F6Ddgqi/8
g+1PSxDH3cFqosZvNrBXviajDJkeMVxLhia+1JZPwlULrTVEkWWpQWQOXd1hmdQL
94h1/C3v/oqORZfgWeFDJsAoQdA4ObUSfw4HMGKdrF85Vs9ngFRiKbnFQQXWI8PU
JMCC+pVPWWU6xA8QUc4BcCTWSg2LzHkbaaRYqX7A+o4J2bcX0VV9y1uJMkDl0CJM
D+4/4ATLLQQU8MhWZTCLlID5wMumF7+dewDZwk6p0tufEUn9AtifY0tZ2WCVDX7/
JpJF2da6l55AbW3hqKz8Xog57fQscb0WuQrB3nrTqPcX1POu1y3RBAdzM2DOCsHs
Pm/nrime4v/2EPkB4ZufoH9ybNS1SdFbgFiDzbxhV1XchGkg1JzyT/jAbm3Zl2mt
ZPgg75dxMASRzvbqJZoZTaGdEGR4B5Z/NsuGfOtO7Gx6p09XzDIcafDdjUo8ootw
sYmUP3jRXxd7qXzSejNaQ2apY3pdTrqOvglkM/Eqx6uBW45YcDKdftV0/lMXzy4U
CbnV/w2DW9jC9Ee0pBOPAgftyWoPj60zZaKXv+5wsmQWGyX7YoX1yGRdcoASOVFT
OYQl6DI2YVKUpdnCfoCfRGBo1NKt8tcT7CGh4xx/U63uVTQEGuQcVsunSlvL6zwY
KIrenhTKiiQuJb7r3ln02FB0mso8TBpKw3Nvrne5ykPALaie8bDMjRXUtpdsFWmI
tysof43q9Ubjiy0gQ9udCpRAPXeKIKh0FPw+JMd5peEI9QlzkQLlrNn/Flvgs+Nk
Zf3a3JX1L9jmd52X1XXjzNQiBiEw15GjlgpXaQ3Uo/QrSwU937KZn/j52EZsnVP3
i7Y7Z9WIYjeCIKiam8jeKDpgOw2J8RaHzfZO4witpDHDAZQ8OlHKoweI9XY/Om3z
Nh2Yd6cM4OzGN8EWaYgUaB+aq7fpGPpMezbctbHQ0UvWzYDuDXyRdnNs3ajKeXfc
d9VDL+unNVwnBWFEO4DTbvxcvSNDDy+orUJ3sy9YzjTnO2Q5MRbfJSRu9i9NkY1u
kF6DSG0RavLkyBaVL/NCcijg8q10faiBpBETlUWEwh0UenhcsFS8+XkETYGjDrb8
Vmd9BEsqfvvEWvw8FmCSsmjz1fNdaREEwNQkYzLcV11f7tdQhT+HY1mBFY5BA17O
QbbXvkP+O3RJ1TPbhSCwRpHWGPa/ODRui0ghZvAaFIFrinbAGlS2xA1M9Ww4O1r8
EU49dB+0ZnCCZUvQ3UkVBVNv+V445rSyOiMhCqSUKhb+O6/Ji1JceUM5iJkkND7c
nxtJ0dnfnoBLbGRFJY1qVqByqx/3KhXKWqrILNMwnDgZTxG5ZNHl7CDOwziknod/
yeXnk4uY2NvInF0K9KyHih8r0JWuLsXDTUAZjw6uxRCIjSapNqdcnV12gWLCi2cC
rq5DaoohdKquFODIqa7TZRH93v6Y06ta5GAYl/r/TQqAKddcAS0noi+oJtDVaWz+
Vmq94KwCYNW2A3nX1ct37uQYLwW5kPIsqREyJODRXhXSpgCgPPdEUBwal06VhY3+
QebCfP5urOHI+DKA6WwCiOnbt15h9Z0DubCAdJsCm3HTePE0ayfVop58Tk3rUKCa
tzvtEaqIf6UjU2Rs0cjqsMqKxWbPkL9f7uTNJ1JNqtuzjAwA+ZixrQ0dAAwesZNh
viEu9SJemB5ks+WlYlDSoknQ+MhAZ2aK28OBlNcnHbPWqkg1ejmThnXocCabq+nF
ghvEScE68aLMo2C5y/v8ujibOybP5I8z7ESykDq93RbwlDdfBQ2zXa0/4YZTGkQU
1VJ/Hadgem/auGB58sFZAOzgWj4Aw9k8S5+GKSCbb2XC3UHSwi+ODq3rTOnLUvhT
OFwza6FcdHODhxBQhsTRhWEP5aH18UKIA+Nc6fGIG/G56ZyDuSaNpNvqsiSvs4ln
2IcJe4TgnZ9E3qtBAneDhaRecq3zRk4mSYjWLDIEnlicz/2iHe5KJVqd8eWPWkbx
oJhqo9VH4eT3jdfhKJ0mJTMgUW9gIqegV8S56HUeiBCQKOXl8ju0bDN5gTsJip+9
/QqgL02F5Y35CMQnaFuoesf/aTFLsGhu2Ew9BEqQ+EnIHKsk3A73VQ9yMvLgFIsX
z2ITPftg2m9y7wfnG6q/vmyqqFyuf1l3lVFsqH+Xf1Gsd5VHQWLtWgvXUo7y8Mac
JPSltCruGffMVPBDxlyuSZHZHk46IiLSwDnMe2cQxgObzUIZEsFtVBDkYmhW+Hu3
cSBh0QApzn5oqMWNdlDP8shHKXDaE6UGjI4fhRZvBSjPj37iC2r1jqKXfNviSsW8
X8emsiVhwtsZrRngrhh8MhgoD09SjylXgjKdsa70hzSbUrMEcUpzcNd2La8Cb+Yg
3SL94vcnNOHrSOlwTNIwxf+0pSaKgbb4UeuYCJ7WhYNN7diavAwlLGQiqDSPb5Fs
IAzAvRENRN2ZppgJB3aCcjGe3Zm4pIq7YhdsdabK1YbqI7Onp19QxDwRSfzi2o8v
lYIdDOoWWqYeLxYwDx32vKY1sulDcDyVWrQO/a85dFZwGe0navXUuocCc8d7c6pS
4lL8rZjr8hJJB7kOQtG5eJzKB1lRe0oCu4fqWIVPz5ZhEl1vgWA7A+WZ6JWArdGq
bZepq4aAcw2n3JO+38elzCMccvhVke7ggCJElBCpH79zhu2TiVP8PRRf6VIYWF21
UJiK0z+77uykrqIBMpLXnvQkv6GMGwCoJFBHS/elXIy9Tmdl3BkrVfEZevKrTcEF
JUk9GziMJCow4mP/G5+rmMOwKXQrMjPEwTY9pQx+ktDBVhxSwd5ZAFRznkKIGMgE
mwsFfokrx+7k89uGk6f9EPW1Nm3GYhp95LtXZc06pmAkP47xRLen8ySnXcbuGGjf
XiVLZP7rJfb3P6LM53Dk7Uo6cv/jgTzqY0fVl96k1vBCwIhyvuR5HXWAbJxES068
bkXwxSk8Q18oMDV8nNx5wTPvLpxNQuWP/VUiQdoeyDDlBv3hezkDebCzvaCYP+jZ
PXfMiibb+Su/phO3UrWhQKq1lXK3nOgMGddKCcD4t57wsTNr6/bcXvSSaDKwaKl5
LBUlhSISzzy/e+mAPin5kJ6HPNGdwZ2GX/DboFZaIz4fw6SfaXAVR6ssXKaTU+uu
nAfQeBkwRtcl1oopAVcdVCD9mwBhCtiOTsVrxJ59Q9r7qO1K51Aw/L/806bWUwwC
CrT3awkKDcYWwl+i6J62L8WYmB2dmmvySt0Ldhi570AF7WJrBYC1/AtFIs5ODzdr
odgYekkCOGKBQzNhlYLXZptws08GfaGAeuRK1S8jmgQUZimravE5YUcp6GLrfjwS
xvZtTvMDoVq20YrJMQui2GAggBmWQFJN+t0b9TH25QPIl/uoBa4bkExIksK4FHJn
L2/BpHn58Kn4OZfav8DPh66h9l6PfrDezLhQUfUmpyAnvgPdusxD0ZHWTBRChmTa
G1vBa812Ye4LaQ1HnC5fBjE8iMnClWrmmqJ+twsA93gTzU+nQsAfTX2DgMMNjeK1
1TqPno3eFmoqPO5UGJLrKlbl+slGm2ff0ngbXOuHcNfGm4sG7MxDCRl2uRb6fl5E
7HsD43683MNtc+b/UP22c31r2Rcfc5K0x5uk5LXLJLXMeYOSSF+d2kiF1ES9wyaY
RehhLjemV5V0u7/4olphFFWJfthbA91k9YeMj8zOH/f/LAOluM+t9SlU3R5xLjKV
4e+9etDkKYK2e12+xSnBznLZogK9BXjpnLWhZW+6hq8E8IOlxVrToLVG0F755rmr
3ng1uH29OLiMg6TOpWQSoNsmpQvXCIJm5VdWC/MktjEX76zzEWbRprjQEIb0gn64
hueY83XE9YmEB9AcEDwZQ6IK+MI7RuJO6tcU/7pkliBtBuhrG9J8GGeFLZsbP66L
HUhhlogScLoxshyi2wmHYE5v0R52YIEIlHqAYkvBA6LTKeE7qCPvzF2WrzwS/S4X
rCGidJ+JFXRVSsfI1W6+mUeaznHi1KguIOv1Xym3lcwHwnj1ysNBepxMzhPVuv8j
aR7NMpwyrYnlgwRZuUv4Ozxug9GbMYgkpxkrFwaq6J9KLkuiK5VaKIJoVdA4dlep
q0CJOpsBuMU31ouxi3r6UG+RUHWebDByr1a1GLHruN5Iw4BXNsV6qQs59jAj9V55
3B6nwBvwlKxEEVDWTaJL0AitMRBAbypEYkhiePmMOWveYMVZrU0IZ4Zy/9H+ds6U
XTi96z9JS7DsYG0vRRdTf6en8vOJd+BlUE1LuijsOLiP+PDUDiEt8YRxw5B15cUe
BDg6If+4C2sFxVVqk7f0aN50p3v+wVw++haRsd4hzUy3KdfUtDxDaaC8KYT4oHoN
cdWzTrUA30gN64mENAgywiJUZDdZp2DyEamNHbBW+81RPSdCKpkE9oy8jUtC5gD6
1Vl7XHqJ0x8TTp2u+k9xLIYJonreuPafZCWTD6MnKv53JBk6C2kctv2FKIuQVA8y
ZXExf9GW4482OTYJofEhnMrfTEXGwxxWwqerqaZoAIGbmLT3hIbXg5fNg4DBFTj5
bDSLQdd0kzfj5AHvPQdasNQK1J6RQ2/3GKwk7aKxJe0GJJ8Ki+8YrGxKl4GapO8P
0GFre0nbnvlYJBdIb+dNd/91CgVy1aYhBXG2WvkUQhtJiyRhCiDoXV3UK8xw23HZ
PjeBMIuXkufgqsnLHxXfHoRkGXxdAFDa+4TWyOlLEvQIysTtEzPwVYut6J6f7r26
vjEjDu3OvFOaaFYa02X/9gyQjYgGV1yiQZS097wp38HESm8eWoTDmrfCIRFuRiMf
fu+S2vEk91cg+lmhM6FMxOSwa2pejVj8dNMBoOqZdb/Ia7ylGnY71Qv3M8+pfCfi
0dTmIe3nB6u6STibRzlWqYWI95ie2j1XI+hEX662D9A81p3Gp14FhSnWXhY7WJ5i
yVNClsqlbnZaC8FcGYK29FW5cuYVghk4SrybjKMLhSfjsDZ7KRDM54C+hwy9nCIG
rKgTEQxyl0ZndNPwMoHerJNLsLPHEDtzH/gnGXgZ9+aZax0Bp2271pMB0ukgxj09
9JovYSeGWknOF8oKPBdsV4zUO5DrQlCqjeQlwnSF/K6tUp7yaP1AZtD31kpe8GYO
tb8BI7W/K50EZ0JRXv/LZbsZPoqX6hbwNp2v3AxprGh0qAqd313x6puCnQyLVRGs
ZZRH/nHFSKMdv/h/8ligW+jAPEU3wsTSnPQKgfHvt7p0DZyk6NQbgJvI6eEcKxJ9
IqAYoEcyPYXQEingPxmxzDLnZvrRZt2L8FqBRcTn556SWbqY+QhJGNlGh7lSc67b
8QyJAVdRDCKdfP/OhNsBAyP5m53w5LdaVvK1EsGdVamalFbozX/NyFX/iVS+I3R8
i8tVJGRgQOH/fjVJbIm/91QG3Z4dTtId5ensAfRxq1tTGISK4DJSKwLArfJD1kpW
I/aLG5oo+U7by2zfI083uov4c0SOs6Y/bAPBmMZH1rgK5WWZ8HbjgmbdgUvzt9k9
2CyzsdIN2DX43k9d8ETSb+gyYE7fS859m/fPcmUk3a5cLAYwt8Gr6hokR7m0Cyff
EJ+rHbUEUbwJzKMrbv7wd4rOU6FSKOjp27xNe8s5ZaxdB07harv5hKtR8aPcgPMp
48UiNupYEH2AJB24r5L/+Vf8XjShwuT+W6qPizbRri5GpcYBrztxOQkHKtN8A7e6
85cnHKtzFCJADqVmDaZ/1eEDgeLWqYNLzMy3Cp64/1beUb/EEXSSk/N0gnIjLWTV
3NjCnFv0W5kdm5qEXEvZ8NW9A8xf3uVO4RMAEYHLbiaRgfXFhVq9DSKucAhDKInz
AaJIvWs8TcI0IKuN2QrYQ5egzLWqktjrrGuRZgJvR8Y77iu22y3fpC6ngpZM4+O/
PvCXAAXvWoeAgLiE1yKKsUU/q00K87zN22S78NypCBTwEdyP3xc2oxYiLo6DwRYn
ZR3LqhiEd/bcDRB/15bwlDp+6OM0I21+3tjDRsGBOG/PZ93ybRuduxxJUxZdtvCj
KzJFSsMZgS4OtlkXl4PoVtVagkz8lMVaamiTIatK0zLFhAX8KdCJuoGO2EyMXZzV
Gv2UjePpbrWZLG9O6+j4TWcSy5G0FDavtli5k+Lk63eJIyGXRB0LlqdOBcb1qkOL
eCQILPQhILGRpoVJ5gdm+a0iTEP5S0DLnntNW9Km/ueEwAnLLRm7NXpySJcweSrc
Nyi0zgnY7xitCP46zjK8a9kCJhJmI+9MQP1zgrBqzcjBuhMhMEhwuNYo6Bgop7HJ
NE89yutscJ2VquBtuuJ36mHBlcq5Rf9SHxAwRglFetqI1W5kHi0JCWmxxfpVTQgs
qZpQ/psQeYOGfMbAwOdLmHkxCodYDzP+6jmF/tLbKMxgkbTJIC5X6zxANfZmcAIs
V2pvboff2lJqppmxFLf29dA6Nikha44XJ89XcLLQWv3YrkNItUZr1ZkHd6Ev02tT
x7nAnv0baBH29Pb1ku7JSZ2qs5lsEe2rIQJ69bA12W72ERW8HEc4vmey+AAND06V
1htTLyKQ2e5kCknB1zrpF8HFa9sGeZIPOw/IvK09IwUa3f/wsrIjzlHyVgMD4sz6
O2tWVdpAYI+ck0g7rFfhwwDyOF8uxLYjHlq1K+mYeo+2kp0KYHeuA/5fIOd5fK/j
zwaSjz23W2Hkp7LhmO943hGlU+aMXSmYZ5V+C5M+o5v6uOG/p5RKKYzRUkBmNvyD
n4mkRd4+6mQOtf08+wFOKoMlGlD4MggcX0cum7NuqXV+nbWgr0ipBTPjDWQWilL9
RClT6zA95C5lriys1qiEAfNComjJwhZT5rSArSxxYoJ2ORsEQ51IoU8AQ2RhC7t6
sfdCxSDRpG9zXqWP8N7gGPZXCwvniHx0Bv/gO9M+OA0vMWBYiIizjWp8djV6RlZ8
b0VAs+5i8VXd8sb9F8Ar48QRsvddn8jVWgRomIVm8+gE75h8mqKOuDXnVSoVfucF
3Wr4SCDsiHFgQ+SJQibkmAW1Tq/SReDoNSaeY0EpefExLW6/93GvRTaKMxSCltPl
ATzFIqwOFD8t3T9pk5lr0nROxChS/7HrfzwaSI1KnIfvJmKyes69qsRh9ePFx/hg
FEZE4AZ+YdtItKxT/mXEOPX7C5hP2I0IId+ckArXkxCi4tChnwjdtdhykhmow4IS
ihhTUROl/f4kWYMCP6HNhfAnabS9JEA+MuQVhncLb55yoGjAd5l2QLNKJXMNjEIM
IXvfEhtKbx71y1KslwBR75jRPyr2su7mCGVWhVnsyFMzLwyrZG+ALHhdHhAsfXFo
7ffLeKti7YkucrqbuaGbb0y8wBgJ530L1Lnnhh/g5HLWx9PGU+4IRtSxMfd2QzEM
g47cdq/28VpqV//PJeu48NMXQ1+s+0arusw14TBmIst9VPHNuatd+K2YhfspJTDB
h3yDuJRYVorA0mBmQHcLwsEnuSJuGhzTPUmMaoqFU0EbyfCA4HKmIomm2/eiaJmP
LrY4+89mhnDmwQ7DsjgY/BjFzI3+BqSRjqYXjTvBDqYmn4DMAMJ4v2geUqdqTHcT
IXLTYYvcZ1wZyTDLfSfRnrMy8XJNRfP6Osa6VVmdR6/FdbGn1WU9HYq9A5axFE66
q0irPfFF+VlTU0+1A9fY8zbkSSIBzM66VmWuld/XIcde0CAe5g2ameS5Hyk3Z4pu
uyTpFM08ZQo1wdXp97mQbIs1f7HjwxU8a+JpWBUgoQ88xs2Fl8ecGVnuN1WQlwfs
RQNMs6bX0Z6SQT9F9tCyFL+mJUsD5mh6rXbElAMMKrXCgeyYZjOLult4MK8MBobQ
lhBH7jGW0JDcaEbXzNTi2yOOLhqBtlqLe/J5j34YPOlruQHqX38B+pshlYlOcZ0F
TPVoD5DCr86VHwWZJj7Go7+fDFcco129l9H+TH96DqYwBoKpfqL+kgXlE+hgMVXu
gqYEJx6PwaC5lcNubMcRN+79Krm1t7GJMLGDdn4OgzonQOb7IkRSDkvl1ZoyL6gr
K6iHPHaau6tBIenDD8OrcVWnlu/yP7CBWwvqFmzlPP2TY0suFejrT366Vt+SrMrI
XIBCBFc90CbsWr9kIgJwBGuok3qI6n3tzbZmk9FXITX6mtt1T6r/kqO26uIAjDsV
lFtfXDcH5i/jfzNa+gbq3iGMZ8UJk8Yx3Bcvk6xxfvh44tdho66GByg74XeUSle5
o04nETg0vb0nldRQnZ22D+mE58IRYba5UYR+6i+78i/D4mV6vLnTsTFXEQquHnNh
gcOjFetimolyTLxM/L7VWEfSdeVo5yIHlXbyHUwg5lf+F3VA08YmnTZQFHaPUZzK
17lQtwGpOjqgACpgU4V2EIunFqg3M5BGr6X6ezIJEMzJX+UM7yxNNxUqx/Hl+JoE
8KUsOApYwIVs42FT8ig0grjqpZ4KtlTVlvXS4bDdhSrl/3IjP0qOGkHr96XGHRGD
2jDA4KRq77MJp2VXISdjqhTSjsxuPd2yrlDP7nd/MNi+NTZLPUcbWSlgvg1GQ1dJ
AHvzX2VMwx1lA67Lo8UXs0FwNdMxd4TfYGfCon/n5dEtM/pWiAj8H91RbfHEVNwr
MVyXFNpvznMW26Rox8jLGmUA0hlndNEJsxE61NCcxW0MztP8Kunbc7BhUp5QZbki
nHWXVf9roLVv7/86OW+F0xHDkcJAruf8nm+pKk0RUAA4BE2XtCrPE9hV680KWuBF
qW4FCIGejLnPVH8+1vMF+elAjvdY2ZErsR7bBXeqTAhpUoM0zC3+M/xRjJkwd00J
PfKCWAPW13o4ME4mOuKWOdRzbDK4adBi6eUt2a/PhXQZM1vChN0xrP88iU3ENeIU
UaWFHLAnYLixNS0UNBvNdPM2sbqW71rG+VVbjgSMkENAkoPDZ2pRcgDlrc1JdL/l
kcSkS4q3pyG6olMuGFq70CYfsNik5sqF95WlTn/+IqeHXXHxZZJ9N6Tc/H9zu42q
Ac7H41aRQsc/jeq6UPS+nfpXFShcfZUQd8fHesiSc2hyn2vvTkmLSeGarnzJ3B0o
ASG+N2/R1c/cAAU5wIV0R94F2JTBFzRf7t/xNGvz7KnXoaEWZHTHGJcU9pZHy/C2
uxEEbkWafVRnz6kELR/fUxKvM6hDPtpGXlR9pl1qAMgYHV8I93yfpayrltqmpCK/
SaiGKD44YHgSrp1j0t5NpDFInrohPG3rCXv3bpNxlFGC1BooppLeXQXej5rowlrJ
k2GgCzualy60r+F/seJrOu7gJmlaHuNB9dzMZdF2bgUY1mYt1/DwYmzo+Oxquiys
z+sdCb4WmjmrYM/ltEkZ95pHcEezoG890Ij/vB8uQdqIROqHxTLSCya31Od/UPox
IdTukrZeIHEz4TviYvhn+skuvOO3EOtQXou27oPIysUe9ayTMf43xCGYLyKJ8R7d
SCuA41TvD3WpF1GHwJVZVXMTNllhqi8lZrq5sKDYgHCw37B6XZCk0Mb0vjYD4gmS
+TlSA9W/Dk/CfsS2ZDRRC1pNTQOFzg0DopUk/kSi4WPji6Fz8PEniv/g8p7x2lmh
g1HrHHheIRGTM5NDo3MAP02+SFSyiaVd0AMdVm2R88eoNaRS922EEXfZSpUyky6V
nWtgV9C9D7JAv6teI5uCGHmTs94YhNVSllanGGV1Pvdg0jSxiq6xYzKR14kQ1oqy
mNKQXkOqZ8hUczR2OAiKDLgf4FYHkfmaOffGKs0rypswIKsYyIFlDPbrIha5dw7P
stgdO3lAgFg6jcKAktq+fFawQXMFAPkldqc5xM4zmESIJ2wjXd9YPWJD39jkuAWJ
XkugB2NR6RjOPdwuj8dZv0D8K+d39p1XiD7ligVpcXKBmBcgpB8uz+dTlgEbK81J
mpTdtZReRMvvTdbNg4OmWETp8c6atOFL9LXOIiUvXHWDbFvJ515DfdD4sYhTX9e5
oiNliWRNtgm5LjmRNBfwoaM8ULK5gJ8hBTpYVIAw5HZjWhrZ8x35ofvrW5gjF3za
e3J3eQ7ovh2CqgMFJeJwjlBtDBFZcVNV0iFGXDw8lUCE8fHj7ttrGH9oi0qsFKnG
whU6XAQ0i+aQPCzIrzImNMF+JLNxHgHYHeKXRjFEDK7BuQ/yCR0nCfc/GGjzVPz8
IVMBFxs90DPPCx3fOddJW8n2xRHZ8RM2cqd9JEJjBNbMdeqtA7rZGwSe3ARdCEkf
W9oooh5+U8EQ50LL5fh5MRtIRwDs8/HUaJXKu3/pdX9aqZHZXkHgZffizhBLUvG9
I6tXVCCqcivAYds44HdtpjinYa8AKJBZrdYJe4gEd7VizWyTrVbTJixeb8tEL4Fs
/szGhSVKSp9b6BJYHzmy998VlrBlAg9f1BrTEyexHtuNM7/J0oyolFKS5eCR3bO4
ILf5GipCCAwOs+blmRDE/EunsTd51HhRK1N7Md9QeFr7HT1EyY3GH9qBakZQUnGz
IUT20ymWPaU2I3X/igdsOiKi+macVztnb/19eFOVBiwLWuRlz9FTOxcb1eJMPiZr
5jI1K8dQSI+6eo0CiD6XIis2mQFHt8Q8vzypUEKnicPKug8jWQPvSdkDmfhkYnmH
iWKoaH2MR+XmY3Y5J1EfjiKGPqvM/waE6T+kEQkfl6eDFXDpvvODrlbvjB4EVXb5
NUk3ORg/u26boDs6NMZFoe+6Jdj30fU4TrZW/w45C/0PImoRVCAfDqjmxUsVQYXo
2qZPbsmOHJ+4axXEG+1rCFEVIa2nNvhbt/HdkBShoOFc+mSBdG9AVjKhWRixC3MI
vSTz71G+5rgF5LI1CTs8IZl4ZpChaPGYPERDgjK3MBUNa3mW8z/twBcZt3MRlXXD
JNfFVUz33mp1hdFwPRkIAQVARSCraIGp+hT9tP9jBcSq2emSDFfPuvMkw5HMlh9T
u/E4P+jU/eXlzdIBbJCGBYLetZdk5N5zDVIMdVQLZSe7MPIL2Di4xfMUojM7MfnD
gZB3vfVPusZLNYigbat3GrB82UzSv943Nt254Zud0eHV2g9f3hnzebJtK2V5kaf3
bkKbwUBKc68VbmQ3Me9e4fQ7KUuPQY/AP8MZ+aDMJ8A6L3VLGfF5jJDFatSUOAfN
5opNxAkhrFovnPKUJg9eiVWnMW/YmTaC37Ylmy0RCks3V3yCwyz3OZ+8E9wKQz8Z
dxF7LC6IyTTtzuNddbiDPnwZ3c+7cUa6huqRNKPEGy92ZCvQ/wJMEgBb7g/Caec3
aKdFwDTwZhkSSSjxIN7A1UUQCec0x7Pv7+JXu83KW3lmblCwUtzr/kkcwYiI1mXT
Y5N8rOLPtNynDV4Ozu2kq8Zpk674nRBShKVbd7YOtUl16GNlZMf0e1Wat5uCzc+g
guugkYBbKlUcIWO1VSYYarVA5LhivC8EdnKjwnUK4+HW5aU9m5+BGctbU2w/vBNp
XoShOeKgCiCUI08hohWxH/br8AWXEZmjOaRZkbzZie1iU4rKRy7odQsx21vf0JnU
+WwiS/Km+ldCGsJmeX/dX2hEPkOb8GUUovvDVikY0I0luoV6xtGRnsxXS7+YBfxb
LFUTiwos2Rgl17nqW5P/mpcaq85y8j2Mmy9/la+cL9TwfSJ6BQLcUFdsIXoFpns0
k2FboWDtBghwmyqbx2Hrefz5niNbZFfZsgnACE4c715sSVZeR3ipw7MvS6wonHPU
at4VTbUtG/fulp7wGMEnpDhctGKs3FaTlbmkZFz8HbIfnbMK19JVmg8mUSufHeLV
ShmBQNuI6huKDExehm642hNUDkPBMfTUfH/ei+ysp68tFeFKhKCDtWk/I8L1MvMC
U7wIfmhRDZxZZWU3dX6yYbrFJtVO0B5FuKXT+VXgNMXPI0Wth62/7X6uAfS7LlTB
XCYHN+bbqr94RjZHzHYcq3vsJcsWmObSvUA4chiNS7WoGk1mlfzz5OozaA46bi9W
l5lJv9lij4fT46483fjhIerA99RsyCh0tiNDnahTJNy3+0Jt4PQQ2r1ViV8u0tEE
gKeeiN+UZKi5m9XBRkWon04WtyMYQZ5Nusn7ao4mIrwSiXebDp70OxmcSnpngmcx
/lmjUX6NGqojUF+Y5pOkoEk9L/pqrwfUHsqHHyGr8WnvGk2wJ3NT24GmEkvkIXgb
65A/DbQvNDrjGg6ZjV7GKhcPMCpLzWCMp7qCcLQgqpJH7VCaldoGRk6cLhPHU6er
y/oon/9L2UO7jDvNjLxF1y/GpaxTtf4u2f4NkCa5+9aCBdvsjG8V3DiQqHpzvMRO
2Z/B83CmRFIU/eK+F+BZcRdE0Xke/BplEF6OKaQqPDkbknaGmbzfc0qt54oEsT6V
CFCe7x7BmfC1QODEw6tCYoIIV2cpqY/uOVrISAvMWwu6LCuaFb7ABl3yJDki2j8w
6nKL2sP+amFLlrKisTlulyG3tOYSKky0aEyfecT267qbiFY4HAvknCwkGJWxRzz8
3vjr5HyNHplNw8dF3NJk1eODA2glpjZv94oqsGXskYC9iwsaaQgtRFaCYjJto+wB
5U7iyDFL3XhL+HzDVpjo5d9Fy+8CJM29f7Mgm6cRAn21pVf3T5ftW60KHSdAqRkE
SeuD1in6NNAbC8xwH9vsi9jW9X03KLZYGYVX4ies7ipvMgTlHE4GuDKbzqg2mWf/
L1/uvxIDsSeah0rsZ9JMXesubdPfT90MuF2yorWqusrbnYxyDTdJNxnpXJQUeMUz
4EXzg/lXxPOZ9xjQEHXn6IeAMx1jzNIimvr/AUj1cgzM58pTxKhiW1bencCH3alZ
t0R9mfKu+6fR3tuJxj2ru9eXTxehGyJxmfye9cO7s/pVwKfbMfpLpFytCcZbowno
lXxoiIyLCF8Cswr82SI3ixvhk2KYYfEioJghWXnQSDq1DDUPpkdUPBOlZ0O0TnhL
M4Ai/0LTfx1z+T8cqzz4IqjM51xs+VS4U4mGB5IcYUfHuUJ6xScXi5UsoVqNbXTS
3BvNWXMKfPcBp+4TbRVOTjISF17Sk4CGpG1+EcoJADfoDUWWjyDCL/dUq9tHmpsy
CItnM/fW7chuYFPt2dCW+jxVNMbClzUbfWie3vNbfcMEbLZYn17Ujzex+M9OIS8x
0fXzTdkentxvxp0wCxDHEAfE5rcQLOt6tqq0yhgcFk17BJQMRoGseHW6vewBOF93
xBrK4KMOvj+si1wiEhopX4SoO6ewEsMzsAH/WNlz+cwDOSTmttRlxNG4jx+Fb4Ha
ZOxdGg390T9ur1dF6uCBgGiCAxXx17xMHN52rPlYpK4Y0oSY5XIfDHNkWxHTxvHU
cK1tOuuiaZULMVHq0zmgGiT1tqr0JwrTYvR/8JClh386O0YWMf7MjroRyLxQmLxy
+nU0ZvAPeDiVMt6III1zIRcholK1cXfwBo2+CAzRiXMJWG4Rjuv11Sbu83FhMkq1
NxqdrjjymtjSXrGm9CcX9TkjnhOlWS7w7Sk8gDQbUYG4v7ldGVjQT0pe88wyQhFi
xaNdNrkX61A1MACicGfX2BLt/j1rmJ+2muWgJKXENexSujd0JEgz6kFEzltYe2K7
tcfezftNeNOK3VVDYdXwvgf7ZUdK7LCYAJDmBA8+655csEi19o3G2Z0kjGJLJJpr
jqaoT1c3l4FZRYxsij0BSzMU+Mr9jt3212iIFTMFWVhpOrvxguvzWEEo+2LVr+Cl
74fnF9labpfyzbVGqfi03sqQ3KGHfwgJDQ+7Z0Yq4WBp6cXzJW7KvdyAFH4bqIm3
eSG/Q6zGSisbSzSDwdWffqqojoYyl/WB80P25BGEJvprP9tNaTGh66OEaLTJFAtW
d3/ZYrjntwyZ/JJvkNwDVbzjSyr0pa2QDY2KJSMkhZZhtMyZJvKgYxdwQTpJyXJI
8BN2024kMuDbdMsbnpWarfvRKKJ3AB4swAiiyiIBCHH58hWqRosU/1dILWqzW32P
lFiOMXEAtkC5PJDFpLnMwO+EnWYD7n6JMm8z63TinViyHspgEmVVMZe2Nr5BYUTd
yv0H34BJ6F2O/RYcMvCBDu5k3rzvekVYM4R8pIB5XD6UQP258YSzG9XNgeGdCkDT
ejS5K110THVyqosI3k9Z2P1hViqn+KlnEfauZjZ1frUDF00WYQg75ZsONQW1cKOR
Ge6vMUIPXgvORr6QPYCsM1BVMUh2lgg+jRWcSj3+sldICGhlRXEfPD4H2HmbcM/D
pAV1PVANN+/OesD4DXGJzoEC+HCrGQ3kzu4yA6ZcLwCYyvj3CJydOqnaZ+aIKcWi
BR3jZTukz/75af576L2JLBUjOYggaU/kyvG+9QbhlTQtruhIv+0WwrDhEIY429+P
FRaL5S5ufoI9T9yu+5ulfUxYFkVn3Z1X2mf04qdhGuoTeY3K4LjaaJsEzHilKIe+
oFC13qi20V8RE3e5XQ5OpLkJI6AbvbEikcMbvXR9M5yE+51FNY6CX0yvYUm0nV9N
mOsxA1C7XpIRkRAVs/vLDL+ajotC/BHTDdkGQMPn6UQLHMgUfdFqx0KNdJGx4nrh
8OW2pMmbrkb9lFPrVnTcHLxju3B9wOYrRquy/78ZkcUFE8s/tOIJz7XX4FjgNOyk
y/LB3AC4tqQwq9UGXS981W+gElsfcSzdX6PTEOxvIihbHIKvadKbOHzx6CNZls1r
knZR+nmrVRqoWuJzIP5NGK6g2H17vNXNJd2bw6AGWuAgjmSrOIN0Ds5wleGVYwvv
PnLg7KyAPYyuQp4tJPjS90YxCQk9zbs31tX6vToZvhsoJxBoAxEXuixvrmKeswtB
EwtTwVG13oKA0f96aHaZuAwmXy0f2S+FbVdqgn42YMnLmkcuzmX9qDs2qZS5yMWt
iG3jGSQRY7wAKYUUcR5KPd7XNAuOhmDxNaLa7JUg+vsOLvqynD6GDSxQGP9hTctw
RShqSSaHh36gir2QG7xbqenIQnxbdvVxzztIBPaHI/5z+EPufwatjl5eZ40LNtE5
UjH7GvoeGJHG02CA/D25epaNSV4tZwZtW+IcnYJDhCp4SefE4XGCS18KH1sPM+D5
SzDjnkDO9ucamsYMzsr4KnT1uYWmF73amJpJ3uKlu2XqkbuEQCWee6CR78mmJ0wm
KtPJkcalc9xKCZqNh/yH5cvgagsQDEBdfFQu6Ct9GzvE+9ah9cwh9AawRfSWxUUq
0Q84dUyaavYCsBoQ2W8dJr20xXVPw+rl2azhyydKRp9lcdeFtsCNtEFQJHcAfW5v
cYUdKfs7OSjn9Ax+nZXJprRdVuZDmYDtQNw0sAHrZ8e45wbOm8SC+pC95FEdyo1m
szXLe2sE5kL8NkA4W9Aaefb8aATp478FKM4CwJy/o5XL5pJlO4fPuxskUrkMnpkJ
hb0EP7Fquis0m3ciAuY16RbM52jkk2kSEFfr01Gw+oo86YqM9lhW7snVC9DzVsGB
oF7nL+a2YrahdVMRaals7qQtFrYn6k3NFE73nLwoV/7VefXXWJr4dbjK53ukJaDE
/wggukQOPGv0SqDX17uwPJtYcoYx6KrcCaNjItBuxsyK59qYUQVFgARBVAHkgZWx
CGOqv4UKn5auzWX7BOo66X119qdLbHob/OflL4h+wf1x3jbPJMdr+rZqsIihYtqp
7HSMzxm094hSCvJN7aT233qzHVdjYJDo59uVEMo97M1yMcE22epWB+PffoVyN/ky
E2T+40/ybgQ5ILzNtmC50doWa7A5ViMpEGltnwubp3oqb/0zAvnjQ8OfnnXlMBzI
UOXTnvJvVcMOgoeQZ3n3vfyRrwMVQXPKOzJG56zra67vGmOLe4X694R2o4s9wXQP
tpgGeD1xQUF5f0K1eyvdY17nErymG/OKKhvNlsVGzgwMAUw4YP4kNRJmQ0h1VFWX
AAorH64HcHa96BUdDUiiZhuqr5+OvpQ6+xUAW46W3kE8AiTqxQudq3CrUM5yMffN
u9rhlHfWeSDzZkcxniKuAMrkaKN0nix9S5hNCDUueNwfVagM7Nsuikx8AezabDgt
EBZHkhie6oHZ2zutlonztA/HeJOJxqEwoX0xkRcFuoWyZAWlj0dMiwrA/T2HzRJX
QR8x6x5rl1io+U8VvuRvQUgKumsaxUouzGE8jeqcWEL+RYSEI+sO/gnHuFLgzOe3
sjFRsmlJOhWe9kqQgE58PoS534JKp19qeZf0sCiC7xA8AZYwAZDGX37oqmYwcp+m
cIs4AZOvXzmtOZCdNbe65uwv6Zvje5Af6jLy8BTsUP1jbn/LVPvLBtx69LrijpzI
eL8CvxIjvOrG78DKRgVQEHHHWlyJkrBmZAMpy2yDVfYqncqTTufxiEGfZaWSnmzl
51DsBPMip7YRVA7iymxozn2SMC5gp6Mpsk3+BkqaUrAuRqGihMADBO2WQRSatuRP
nuzwN1Ra63whgUHwyNUZ976qvGaibia226wfyP8+8L0mfykQcO9DkLerO11oRdG2
nwLXyQIf1FWjtWxx6H4SzudjlrDqU8tK730Yb1ZDtlnUM6gz325xOtCjILKZeEWY
Bm0rMvod8Op1s6+WwNJ8Dc/QEhQW6zpQaOSNjGOWPNtWf4tJJwDo1HSVGkbsXas6
zKprO/qkWZLGMoh+847tCohY0fpQotLhd9HUqhvAbUKdmhCuFeCq8NvCl5N4DGR8
nWM2pCgdLTp6mAAcJBmAxv3DHULjFrVeh6XCdi8lRZHsPRye5kUdNGGcP4S/U+6p
JNthdo8cTZ0MU4gCerVWNPLtuTWY7TBiGkEovIr5a6ktxwLr7AM9MCRuQrbvZ7iI
bkb8l/I+/D/eNpcvRDg/I3C5rK/WeEZIvwSiofENAJCQ+fIcgVWRQbF5Gv8dBfj5
9vUIkepYMYqQI0c36tOWSR333aTBGXaqBny9XiZZZ1io+eWp87yGzNRGNZtjh4B8
b5OW/aVG68nKlDZz6mU0fpAEBlck8v1uBT/QOkLUmuUbGC8WqwMRuEscRe1yxV4Y
UFSDRDH52y1QpNhXx+qW/sFfaFJ+LhWGXYtzngX1gIufLHGUCPSVOnWuqej4t23m
zDwXB4fYLMmA4QI9o7DMxpuNFbVx8eZS5c9CDOTwg4bEqsZ03/qZviT93AtkK36p
qPX3LRirWBNORbdEmqH4CePhSUIisLlEKJ6vD/3uz36jjT4X3obbaiY0KssSCMNe
Wj72xr775qlZoUkU8YKx9PhD0Zwgr73R2oMTF8N2IReAtXNVhj0YGGgIkNboIPH8
Kmnwh1ZcQq7Ev4PwQDBGtrJbc/aB1pw4f5yPF/1ht0UW1hXo6pIGFQ1hquJjLf/q
716kEm8BK9LhPCqmA3dpaiEftza1gd6iFB/jSKAI6d6bWJcT+Z31RKnlKcOL5zce
uvo2Vr1HzKVeVCTELDbif7k7Nu3wJTIvq4jO1fpoLjttEVeRu2ZqSc/fCTELmctQ
eS1Bum+tzd6TXIsHIdJtJuk+WWQdNxWpi+FYkrXLZWErFR/u8lQ/GK+i4LhM1Qx4
2veMqOgeQ1Wu2Ql0kNBAKeoiRhHJmRwHhK/vO0iyZUVw+w0zVR7ofXQKWTIaP5M8
tzrUj0NjQ2IrtZkH21wt17QZrU3xXypNdMVSbo/wjuojv67O2ZwNNPdx7fQ9lOf3
mJQY19omTQ6Yr25uAgRPEAdfVg5p3PGIX1PaB69W5jj1GbKljgPge/rD3Lsb+dVv
UinbRMChp7SIY7jrto99Gxo4B1HACfGDDvpPpoGZ8OPBBAEoGTdwaw9a3iaG3AXT
E+rsM8Woj6SHOeKHv153cFOu8FddJBZJ1psLPh6eWCfHKsXMikZwCtt6+gHD8+yb
u+AgN3Mw8p5V/BDoY1uEaQref01y/nS22Vtj65/5d+olX34FMAEAmGnuRj/vaDl5
CVYEACpHGO14LvoNZUrKYAVzEEydFVIzelv5NskF5YojcOZGN2/pK/bmqxVXN0Gc
SsoNRO14VcIkPvvUO5Qs/sk7zWX1uxC9PFO9FjKtflxLVCiLpJMwUDKKcm6HFXr+
k9GTcRyOrphgl7tK5rA/wLtKZWJ5sj8Krd4Log7DSACOseSx/laGqtPEFKtN+lC7
uIrpf/JmZ3aC63+DNMEKsgKVicopzykQoKdZC9q6S3ZCPmu//sdtKnbFLU6sQ60M
RvygA6/C6rrmDyOVsqlicZd4CVim1CsLhehzJdET1icYBGfxe/M/zXs2icRd2udg
HaSgGPbl+7SQiMf4gLTKYCH+nv5P0bM43/tvrvQmKoOOwQCPk0FWFEvsrstHQBfK
4apHD7pRoWNsI6vW7tlb1Zp1mySr8dFF3Qwl9CVFmykS7wSgH8ffFeaF67W4EdU/
83e3UfvgnCItP56HIkyiFKl8eFy33CJMQIpNPwTBMnxehaN2dqDDz4bvR+QWyqdQ
j9Skt4N6SjuE/nrupJoZuzDFCyDhD8DvqdNNJYl5s1QONZzLCer+nWw2IaTzcamK
m0jPDV3ZCVg8OVhU7B0BrYdPBt+yFlrnOXvZbyZA27n+vUHV6uyv6Mn4Qnvxen7r
lQWl6bKp5uYtFbK5ufQ9Bnp+fWgj7eQoaPSDho3H4laZiy4XA1Ux4rEDLkxM/mKy
RlSququXINfSTp4wmlTlMP2msMlhrvlnqQTjJIhrqNjVgZeaKRvBWi5QRBUkuqnY
+RGfz5KBTukHppOreFHne4DaYr+1Gg6yRyqkRhKt6iqfkwq0vWfbGkIrQ5zM1t9g
VEKp7OQY+T3tSsF3YIwJbPk4NQS8uoa9hUIPtuWWuakZqLTJmcVgWYZy8hqkyNP6
HUgpofSrRjwpMHRLFjSaLDo3hsM9w1/XQCF97Bbo92OcJOFvOlQ9hHfpLXB4FKg9
FOD0/aJPgAbRAUFKMX05NBau+uZB4kwh727Eq74MMPCpm6PsbWWEvQlLB66C0NrH
MGOhIe+GM1bmZuPoAJy9bv00YEyVkyfwSCcEeur+bMG6rSGczQelxil/Am/QzdLR
UWxbSyihDk2xzTpk5otxA8plflDhbTbtbchgNV7F7qnEintKtnC3FwnGz2tcHz87
WhUnBGG1jXNMUI5UEVLwCCw4IMfkGQnDX6Gr4cVFsOHVSftY3NTaG+xJ5AX3e9Zj
SaZ1AaC1LHyhvLq3nu5xtcsrmen9BpXY4a2R0kjIVsTlrLJWSdfIhrusgwNe96Gu
CDndDIARVwZuVTLAaA5rJIfL4oEBAtDS2GbOi4mh9QNkgn3DnnURTf8/FkmiI1fw
SRUUvAspn50ycain+0NKWfcAR9ifOEuFKhRw3k4u+FbsMvXYwwcujPo1hadU3EG9
aK+RMPCv74LpFWYnQaB7nhKbuQipsfs7huWSGG5QAqVmTkXJQmL3h6ALjQSQ8e+p
TotZOoucfPlJs9suuFz48UxYiwj1/+92MT5crRzVElIJu4PeVfnbyPfNI3no0jZM
pyALINTmKZJwPOFGqQku12mFTPdB6zdqgGJW6lrTNah4ovw+j4iTd6Fqi0P7rs59
VTTOXWxkaIaMbMABkJc2XVKdwSg3UvLMzlQK9eyWt48bpaaUs4CCdyZkvFnHwxLs
d6P577Zn1WdlPsbb7HLf1jLEEb0TdUwylCNSxSuj0sjdz7fBjn7q0HQBFR3YWK5P
Cr06gNx+EaheYfJgq308BWT7J8sOEJ9fQtwp9rcN4ivZxGag3nZ5UJfHaSXnSOjx
gfgeaEvNXFB9IgaIGFl0ZUHVOZNHiXGeqzqkdUwC8jjkCdLxbVWOiWYz6QU22zRs
CTLrRkjZFGOIgUAxpRS6j9g4ensz5Ovuu9dvo+7rTW8t8pEJZyQO/fchIcpDPWHj
+GoR8NZzr8dLGMSNmkK78pEI2EtjeuP9c02DbVOrxP9Tel10yj0BXkkhknECvm2N
1c3svfw7q1c4V+BJW4oEtyDLL+bEpJWsMFjqNZfL7SEqfcTu+mUHNNq2Ayxm7ZrQ
7ys9GTrkLJkLdXt32zycHBD7RhElOvdEkgY/FOKzb6SQJspLdGhl0sEd7BRjFh1r
mfcJOBAP3F+aJIFlMfzH10JgoqX0PZ3LIV5Hwogszj0FGc3MAkIRmDi7fCLNbJ3p
IS571YDIAQKQm+YCSQfTU/sLWYr01B86cx3Ur1V1A8HODez4fOPO+pgJ/NkMAOKr
44iUWlI6FRu63pQiIru/yixNQw8RWVK/+XrIe9t19DewTWPSU946h2SbBFDcbvtD
xbbs+msEeVS9fXHla/fV9P/AVJNqemLl0yujiVATvzl5Fqbz6B12TTtZPO2ABNBe
7Qc4bg1c4uDuf+B2B3VTbypcUCGfqQW41D4XD6NSp8XnQ0tkkK7H6mBwKNPlsBcq
CtTApzOYvd9+a13IwiRTz0V5EP6tXCfMJ5HEUGTRgZBjxoVMw8RvRoXSMiEACoDt
Dlo80tA7BRELEr1A/czSYdzgH1F5f+oLkbYQNj8j14NMBLsonN6xxwlQGiMACmT/
BdDsfrVk2ezCgqJ/dvlRwNjVmTEHMxpOyunr+/Go9xkLdRfOGg/HtDfiangB0xPF
ihd9lAIAMZxN29/jUg1FRWT78QpQS+pMFO78jZmBA7Fkxxx6ekW4gMD4nt7Q/Tzd
lmHmka9mJBdaQLOfQnUpyk8HRqXhesMGdowWMZdHZWmSPDyBB/74/L0GtCUFHAyh
+MsFfmwRHTVDF5qP7yLrtdN/NWUqZ/lL+EvWrHpUZUK6rK2L0k0unu9SVujP/TFG
E05jPZfR1/XoriFmS2C2oziGUK9AXj19iE/F5kTu0tGWPClMnDM4cb8Vz96f9VvY
0NWpdHA5Fk5AyUZMYM8cXbzbz7oYCDkXCiuWGFoFTwiitJ+59kgkGWtQPpDQ1QD4
wUIDS0z9QGeyoTObj29IFEYmOQ8556x/3ZHcy1vPeSbs2IptQWVOOiTwfyoMNHvK
EIo6MT47QyazqjxL9FbW5pj2SIcw1mlNg8MqQIw80Ye+qyB8QGoC3CzVQ9cxPKuW
JknHKF5VXk8rp7wLAy/pml0gcUER3/7hKUp7dx8hwwIIQ6DvSTlpFvoaoqCX+r87
p59qCLTdVlN9D+JcgU6Mcw6ExzUw8XV2vD2YHGws/CmLeky+TO/kLYR5b0zujlWZ
7oxaBjvoQJO0fsmQjPc+Anhb+K+UoMmSeCGZUyUqH0T4n1xES56B+1eNjPbrug3T
M3n/ZENo3IqZ/bQTZmynNNPo2ty0I3nQGT9+0yR6sJG3nvbY9fjI8gGkzDx1D996
x6A6AiDhia7+aEdtVDJ2KqEfefltkhPGOh+/6edRrpwSysmuy8Rt9TScs6BzzbeJ
/YcCgMAtICh4pir832i0JJS3RfeoXcS3MkmYL1A6huWtrNRhkHySu+J4s2jUvWXK
rm94OboXU6N7U3hlBcRbr2qISkWChYm7XfKxTrIeAo1hp+POintR073vAMseGdYr
d3nBssVLDPzv6Jc1iH7MEaFFzWyq+r3xC7Nssbpf/y/DmfXhG5xG8MH+v063ZeYO
InBHkiWyb1VvXIBHuR6T820HqahcXqxOOuylSCsJOcJQMMYAadPLAqLwKzeePItQ
brzKcuAAJz5zmgbGPDl2eaTrgWtZSXZcr3KRZIg5udNEUrutQf5gJTIEzVSiZwQH
x8+DsLGv24JQkhm4LKPRLq2SvEKZudfyembmKu59/cRtwA1hlffWklXHzn8V0ga1
AhKX3zaaiCkfMbEVJCu/IYbwlzEhAqcXzL+MDe0sXEbCyIQbyXFSgTf7BREBbZ/h
Gl/gsJWlgj0ifsT4Anih3QHOs1PaaCQt6VgYTmfmK8p1NNs/ggZ4usrfxmxmDog3
d7yTzsGwamqHASv0VJ8EG8QePPNug+gOEAam1/qVKKSIKQIERmg92IVr9iAL3xU9
rrM2f/gzNBpQNJvbgGK+1ekWgbRdx2OPKQIDlJsfVw7paBJSFhX8BKihHRPHRgiM
7CboiTV4jEj+R4Nun8qo9Dx+wsX9UrYf+2Z6E8/x30YmNwDhCEwSE4rZqejWbzHn
YKta+TESgXt1C5ShQTGs1tAinbfp211zeUd9kFRGwYpf4Ix66/gLTafpda5UZUS6
qLx0wfog/TNy/9BwUO9MIaLDm7t3HCkEyhxQi2uChWaF2NU3S4AqRUVRrtXPDO5D
PCWG9yb5+hRPslFWEIwpdcVuuB3OEfqkgxBaZ6d8G0m8Xi2Fxj9jL0CslvzDNk2j
S7f5fg1knPpy9lHbvD88/Ffmh/2y1NN0gbUnJ6twl5O4ibLcbqJgd2yOHM99sSs1
kHPe/NlvbDUd/x+nOQWpdJM4ZhCji0zxOtJHyPIeZB8VxQcNeMjXsr37es+m0W2H
XdSLDg+Jzfq2kpI3vIZcQfiEgoyacv7beo/MkPxgg4Z2MmLWaGfb+3VY04c4vL0E
BA+14SJwCzHeRxCgIN18rb/SzcKOnFGvZwOLcCHn+hyj60/uLHYGAwM9bIWvnDza
iTs/nYHJS3BBYoIhgJTIKFbd+uhbYmQrKbRnJgakLeq7ZtTGvYUakvpyakQLzydQ
YF356fBhOUaL6z4U693Hjis5/My7zbjOU23jfAC6dPbT/aswe6jPcDMlrBtqru5t
x+VdYA9L9cnpx9nzC8uyjNtZYX/ok9eOGcof2r/ciguhlTPN569PeIlQ6qbTDvcC
vFbRQ4iYsa0qibaR/V0YMx51aRHxpdXCKbGhHXjKmmYIZH2acJ0p4b62OVfQjveL
4lDyT1c1jydZkXbNM7kcOCcKJT0t/IFIerhxREt/VtNi4BWaZki+uTMxZGjOB6Wg
hRaPpFd39rgy3J2kOrzkDAtmtuAU72//mu0ExvP+DZFdCuJ7FKMqWW/2vw+Aionj
GliQmpfIZP3IpaSPNwZM/JqwdcroaSScXXC1ULF6wK0pxZk/swtPBbgAsVClP+Yh
PToeCnqr8YIHVyWsTotS8GaqXoC0Jw6yk8dui7qRw4C1hGWR6BDDTUmXa+Zwaish
fV2jFQpUAGDnHUXVJzbutDVvM3OX/QwVSuha+um9BykylMDMixxUqpq7yWvtTIvS
NPO8W6/m8BFc/dEW1HTuhGdjD1oo5MDISNeTWlrfHmJJbtU1yC39wUc50ykn4JH3
0u635q9m8nueWVligPWLfbxxVtAqHs1Hk0m3EirzhvgiprVe9zKWmwSRmVgM2h58
tiQxKlLrRzYShDsPKSQDfeDOCYF8THcfZOodG/00k25ijzaec8JbQcnH46LTwWL5
PdrRAN8GLfgvI6L2BX7kLkO3IuHcV2TE+iiZObwwBmuicDOQOxO9EzwGZ7gFjr1l
miLGIvA6IOK5N3/OEQg8+GvJhHp1feA0XnevY1vRGufyyhT69MDfsrbexIpYhVVk
NjDly6HXr1uRPkz5dxGAN1Hk+oxLq5QXg6F4emV1eD0J1M464w2U9kCLRywc47qt
DUB81Ua9dBE6bBA/dOqiJ+RAYVvWLIdhWBtwl+NEcIS1Q2xgM2r9ah2fgDaYV/DL
+nDcaSimhSBHD5C5nxOXIyW29AM1eeMMc2TlU2xUXcVKb8P8kzhNS5twuw9wMlEu
T/NRWCEm2gmpdiDD/gUo9DzYZMed0VrN5gCL4WaNeYAiUy20ShnvmGva5pUe7lm0
/YwyJouk+FHhGCl+Dk1Ixttr9QHwHquIze40BfWHmbLuoAUq70/Zt1/tiOOscyPz
i0W0gnWJAM4XsonqlHDzTFkKX0cKdNhxi+wmYiaVxUnWW8KQsfUKFC+PTs+uElBr
jgT5YWLY55mOGVAY7jzGjpJf19f0f4QtoYCt+HnctbHx8eL3AY1HEfMd56MZAWBe
XuIQns6zbxyIMku0zRGY8IeJyL0gjBFL62ZsLplvwbaT3x0GNcpOSXOey8RITtbh
7bPrVlV3SCunmUeX4Z5VxwXYIf7LyLFpBkqOxDYpplDPvrfLOvo6IgKUknogpvnA
86L3E3ocAziVIhTY1HvneUqZ1LlcGQU0c1ooSEVJQIDQWYbIErBMHU8M54T8GpAm
J9UHO/LNcGYKI5/y4/D3q1AM8CM2zixBSOPHhLb59S2dcewrgxX8QzdXcF6dqp1X
Ln9TYyuJ3YQfMb+mGoF826N8k73594n5ZD1UlTEAZowOBp/aALXZDRThPwqFq6EK
YoEx168hRRGboNDUje7V5cjX3oIjry+Dhk1ZAGDkU3di335lNlk7f1y3gm3dbyGy
xJr57qJB1oWXGwgatfbQ/sBxM+FkOYvBmt4KrRy6TpN5uf7ATWigIA8a3LDXkATJ
I1TqVbkd32kvWli/BroVxsUwM85WQSXph4nO2P9eIXFK2/0BfDN8VzkracpMEH9e
7gI6dwubWWhWIKUeOfmzdcBR3BByf6XHSNB5M8jUfJF1zkvm7VWo73uI/+iaXYGs
N6SHyGul0ySbBHZ6bo9cjO1tiaTY1y2H/PBRDaJejiTopQfHrqMvc6WOWXqjT9wN
iSC/DYICSkli5yJcT3FgIr2SPlBSy42tn1FObtEmrdx5ff5lga8eHdjqRphvuVfR
IUtuOhIC7O97JKvtLejEq99trvew/kvV/0AQpKjxtuxO+AI/XrJx1qGERFS7CxxM
9IOkD1hL/AjpydSSmKFHijJV/lFa1jF+t6UgVRJCPs43EnrDheYBvxzsTPyZjml4
PHNTXlZA8Qp/sTayRrKKOt3N9AOP3JPMT6hluL8oZ675VLI9MzT4+LS76vIwpnvS
m+56wFJJfxS8LQucH4fjj6WAdwlzeIxj7wZXCkYWmhJhaFaqiW+vUlqGOpFXVb42
2Q5I/7ox0uYaYtGrsLXEnGzrItDyT/6QGtOVeZUSN2VdEKHkQseoxwuwzCkVuoqf
AvQCeroJCvv5ievBbgAjCyG4Acl/Lul0CLzpfXW2E+VyUWAwd97Eqf/TM03wOP4k
gqRhgfM1vuOuxZh0qgRWDU27zz06aOf1EoRGpcpVRVzo/VKXlKHY84j40GL3TS5v
km9VxYD4GECfc2H6K/RRPcY8b+QssH7Ix3xn7E4q7ItcV1LF1ThoVIm7Q5pwaKWs
pCnc+c1p/Kb2Q8e4f77/BZLmRPt55+KTOBTgDc+EYso+on2fqBu3+utA9j8tOS0d
ukY6y6MRM5P97FbXFoMkTwQlupCGIzx3JV0hmdSgeBprgAeI1YVgIt229m3rOtjb
K910JBV9hWsfleqeGXCrOQTiAw98YAHM3ooy0qHmqb4M53pkktIRRtICggpUVRsB
RAkzk94HcKqG8VOAIJcIxG95bmdtRtz2Easr+CM4EsTBHBuRygnuBHMPWGuxZDGN
NED2uKpOvnD0qiuKtVL75WZ1R0KRYC5Z7d4KCLcWGAB1x5rciLzp2le/XbsJorbL
0M/kZ+puiImTwR62tQ1eHDcqSX45gbUQtDVCiciz/uchboAGl/LY+Qo2iCP8vT1e
yK+HCFkl+ezZaAF/cynmp3XURkUoox6kXrJ02G4TSlywtQXq3Qj3xfLPkmfR7e6E
ztnlTTRXns3HqUot1XBzhg2w34C1gowJSncC1fxJdEb/fSTfLmhra39jRupxUz6o
N+OUiSM+rtRJWzlSByGOeTWC3wFcQY7DlhFxJWf43a1xcvtpLfPuewdZFxbnVVZ+
CqOnKB7XVBkBrkHAqfQuvVnLAbjLOW2wM4QiPpthPYJxVPPbNHCtrDLCF2fCFQWH
yDeNegqYT3TfExAHaTHHugHuoxcPOKhRNoJVW1tySxhBpwUsRrg7hlZGCLf8Jn4M
3tyxXwoR0ot3JrWowtezT3rtKP2sZgDXywBfSvxttw9yNRxTJ44tKTaiwaaFoAwN
/DYpkFNQV6WliIDf62qldvDu6o6zSwyy3iV96mJePuif7sKkl6WjfYGXFQDhfyEY
Mr8o9xn8V4rF9p5l/DcrNtHhb8/asKgXfNBsjW3nL++vARR7eKuTz/jttWcQ4SUw
P8HIEoHqzLOZj4pNXEh3vs6wiPAweMIAvc15VBLZCZSZIHLNU8YjY4N8ie2/SHm/
6enziRoLazp+smkDpbAXx9FIq/02fWHvxhK3JvhiPdFMWeRd+fHi8K9kNXb5/Nd6
Jr/JTWftiywobwqNgsmnvWd4Pqv7cK3wjXL6CeMC0k2XkSUnzlCWTvVw+R5djIlQ
RbSPKXe2/ggEd8vMYbs9Hl43Cf9US34e4ToVHU6zgd0G8AemLgJbNJrxl7uOAQ/1
18HdJVAmOTZf4yslxMj2r2PqujPxpYWZ9+E0pRqI+quTomgS6Z5fLBBtAZtpdoh3
wACgMHs8vi92QcgmsU+mrErleZQSoGLtYABAlkwVJNFNhAEEHUgsWUExue2xhGNA
Ht37E0vyIxUDvtRbkBpqe4hkJw6vOsfvxEb2N119ZpDbJZqVwjUGInoG5R4+faTI
3xuUmdE8ypj9X4z0R5vfdkkF3mpxogcVIwm7nf15tCjkNZdF/j1g55djwjDrW5/e
sRKnk5sQvMP0wWVvz151sYeT8WLT88RNVBjpzFpsSEAX8Sf4KSjYW8wW4GsTo9Vy
CU4j77WFIe9MTk+EAfuhwaMbjLKqjuq3MH4qZTqhmfXQEFlelW/6OnvTMuhy6rXE
ei5GvL22kNsWEUuAQwm7VQHCQwkCbUw8kwNPc19HSEY87IwC44HlC+qDK3qzg3b2
iKP5E7dM7+x6HjqMoBQaIiSqz+WkurJMU+fIA4BjgYMmIg1qZ1BI5sziOKsciUWY
ex+1p99yvsNw25iMXSUSwwWZIRDTmFzc9dTTryHT6RLNx0FLJBIyqyEmDwJzef+9
UmO+Qg048E2Ffc+Y5weqG0lfritS2GrsnWA9lQsoHV68obyUs0dPKkaT0CHsd0db
UmYAO8J1ZtrDcGg2KH36q1sJWdLQWVCnLqgGNmtKaQlMdaQklk7iauxrwrPR/T+A
XiCPlgijTs0z1wT0Dn0SA57DO326Dx5RztOsWp22IHcnZzImidnq8Xy6/LCffmwS
QHZh1bjySp5SbrcQrpRWRxg59NuLQDCl+1VPGUTI/4cicHNRY6XSK0iPz8UdIS8n
H+diOQ0p1CZpthzHh8uI6QNNV7EdIN+8sm10TAZDSran/pb9Hmm/3GEDA+LbiUzI
KNeuV+2S+5PgQsDVUUHQhbNFgslMKmEThuxj89glBUKSGwlCTxBOGk0uYbZHAqxn
jiniq3Z3phPbczGbgCbLvAEh8osXZvS09XDiLDw2WPloywlNiZbHEL5YupQ7udwg
R0rqEpDkGwylxevewoDq0oN4QyWi1yBfDvp4d0le4CkCCZ2Aij1ELgMDqBnuZkgg
KyuYEgnWjlCSHxVGQ4QG7NVISQ/F0FtjfBl/UFnZUTXpMZh4lrOlHQkdn3W0W63c
0Nier6e5MT/OGNSIH5VIbOgxUtYUP/8LT720xA0FWiUOpPiPILFVQW8xrY861Fph
/QtNX8aY+zmKTa3V1TSsWL4s/F56DTJDS7oIdc1QNoeQCxX8Qzu/KyxOC+lFMqn0
gWaC8gzb6h1aZkeGJNW5Od+vYj6TnGfgjfUKAO3ZwK+ICgTcjze20dLizB7HYhf8
8QaGkfhZVx8AzT9BbTwbw8+/FkGI+t6etrl3GQ9iPlm+4GSknaCKChPJXAeQdwGf
76kJ8vDVIg2xvkbUEc/qH/U0788tkp6zU2gBzHNwPSOjfqcOg/zZSR/lE7CSDsbm
2qJU9OySZaRUHkLIg2VqaiGRfP0JWz+QfVFv6UgY8/ae0xIRC36dSgDJ0R0iA92n
hYS5whcLKEslRt53NkU53HvizsWH/SUrA8BwhyN7r2VrJ+Mwe5Xzy0ueb4eP6MDy
hMERjQoZwAO+NZYoixgq5dm2SXx1Ar9YNDCgDPpsWfd1Hv/pBeMqgtoK1OUyB8nR
fMmphaZNq0L46H+YAC0/GgebNvTWwnYAw70YUdnE0Vuh5plpcbyoxMh3DGAn80dZ
kOAK86a3tF+sYWHJHHGZxlf2nZysAREp0FdGQdM8Jdul7cNbCBm3CEymzvbydu4F
h/9D/dddB0qE+vGvNiGihWK4g2FYl5LhJsxkS2jIyQ4RzG2NTb1L6cqunrPGUuHv
ebqp4JqC4Jg//sZ4FxD6Zn8XzdHc/HJDC3ysx5lRsDcOth2kUhxdvk+wwOP3QLtz
BfnMiAdjdHJ1xj6pg9p4v6I0P5l/fhdAC++NW1Kc0Sd6laXXFiA+/n6MMYwHMLfI
vWQoe4mNhWNbZa1m79EyqDYU8qAQ+7mqYES0coI9j/fB43gkavxugiO4vAFqZkdp
/LbZUR1oKx7p7EU0GZmeLY972anepFoOkW1dnZVk5mryHmNU4hDpJLxKdNcroO+n
0mpDkeCQ8d9ywYC5lQratfJHATmhnhB+jh1sTNPG+JP9KB4PU/5jG2U7J1+Res+L
FX58YAPaSPV95w0P5wmL6nNXOSAwuIzyJufbjIXPodn4rLAZN2NcMc02eb4yxoOe
DoZiCsFA6fw4JDzgGqH0/wGgwayAK6EKAZHPavMmt3gy/Qk3CNn5ofN1SFTUKAtC
bOzHkFIwSbWD/G/rQmxVPRACNk5QX0iFG5p8/P5mLP4Jp1OUEy9wgkxi6vCT4ksr
wOwq2d8RUXrKgxE8mfP+tVhWx2X7HQWsnPD+Efwpz7TeDBw25AsRBDlRDDvf4W/F
XVwoDeCAoRuxBQRTAWlvo8Nky/EG1VsGuc3+KKZcATEojRKpzdWfH+C6jcjoWvFe
N+5xsvXrTXpNKeL+5VlmZvc9smaVZX/I/odSfu2lV0amMFOC00L93jUBowxv0sZ4
Q8MoDwFAFrM+loO51AUSwgEPIyzWKBempFBSIHZEc1Qy50yG4PFjh6wABlbLiPxi
BxnB9lTcEJOpCmCp+/ZoDw/vVmmtaeynAlmHAa4YIg8PsZNW2jG6bfoxzQUz3mze
3qj7mlIorNkzCT6S8kOR/oOyjVfaKDMgyVsLJaG5yhsk0zaRt/wouYmxFIgEMVqG
rCR5wtQ1ZUasFQJwwjGGg8cGmRNsHzTmvif+De2vrtI7Oi2iFRsY9yAzUuKhgBTe
NppVk8hCGNkGFN7OPHN/35TPc6zRx/zVnHCzFlNuU0aIvNnIYqi9DBjFu3t1pZ5x
RiIPgZKDG3FO/UKcx5vRJ8zNFa5tTi97KwgDdlSjIGn3o0n0YtBAb6JrQ6DEOOYB
rOops70iLQ/SwyyHRhKlMAcejAhLk/2UGvZIcdTeoyfhq+/gwuek4c/liyJhltxK
AlgSOaqMVrhTB2Heu+Z3u4rLuWjv+R9+nZ8Fy+YxPGYCVk+B31vTYuOG1q9KObJo
Wz7fqQE7tNCvxplH3uHm2fdSsHUZSYULYRDiDgLQ/QBFnd/yqJyE1qTwvrjaRBOa
F3pYzPg6ftsnVOZI+tjm2hO4vj44opcPhiqvXsGIZLpT1cWKW/z51tEc0ZwUs7JF
DZihZw8/iaFhUCzTkOuSPlJmY0KTQ8Vr5x5WgVnmCk734FBqfAPVOmpPYmyyk8Ee
toIqmFRHu+/dLbAKOrYPo4PXiyecedL1cyR6b2hhsJT004/wiouj29rsVMEZD1Tp
q8ElXjLgB8F4DqhFJQVjh3ejHsG0d1S+vdnJ79fwj0TDlMOQ1H4dvQqoOC9nG+O/
36kcYSWL3tbK4bJA+1xr9g9HOqRLQXXfO8DGBkOZQwwTmDzLqgEL5xjIHcpOZ9Sa
TiJpoCb6RUiWpTijG5lU0FuB8mtAHN+y5AhgL1iEmf5cZlAqt0AaJiF5fSOuj2Dr
XA7HMdy2ApTZQCEuRXOmzORUk8VvdtZMaVcqNY/ou2bOFvG9IdPib0wDssKy+4ya
E/afgfSCE635JM9n/nmZ+vdgMfwOL0BbzIMD6PqrXjrFzA2cR1LK1HZxFnLQK4Co
oze9fXRoTtr5IaTqhIs6Hfx20r2jRak3lcEz48pKysR6BgjN2CZUUHegzobaQSGx
riOxQNrQksa/poJgqkrDxKu+AWKUKCoZDwnFhY0c7GT/oV+00Sro1ghBmenhAolm
CjpP9bWFBqWYiuD381LB2LxmfATQdE0H6gYcjfUpb50D2ZPYkbNdp4vj/sRa0AmP
1p+3kGLhU4f7oQozJcFjL1u7QEw4pnkY68Hvud2mi9/e9+WSgh19bKlLAyiF9fK+
ko1qU1C1OvJcnx+72eBLOrXhxFGCOXu6Cb2ZpG9xcg/5tr7vgikX7FMykptiJhWr
ggDvBcwqjxInJRFbor19D0Pl+AVq1ACEZyPCKiHIrXy1PS53/mZpavjABifK85IB
6ca2M6wrbCfDaEBi/W39d6oWrE1Tx+f9GGV4/pcIvXHVfDoLHkTzasIEnkeHULgS
1RIcYt/8YLrob/2hufmoxo8CZ9FmBpudKwG6T3zED4B+AEM20mTZeIxhHxhe8Ax1
C6Wdjx5dQPVUFLNPcxdcik0DOXF7jpyK8IpXub3QFZopsvuVGPs1s9d0QABSamqa
IpwnxmPevEIP2Mshi2A1wcChAwpiOczyZjK6M3ie5d1kjJOsWEGvOnfRgMovjr28
M/cUybmlzGUrge31do2WU/SptwcR5mlMv8xzSvxZXLC/quYGzZ7WbotheatNKSQh
ts/qqr+oHvRzndh21Wt+9kbqltLDXRBIvhsB923i1xEBDz7SfW2aan1SQmgoYke1
mmvago69MhGRccTpwj0T1e5vKnypIAdW+t7L8tqUQyKMCy5/GIykhN1sMimCiCbP
7C1DmfIsOXydq/BBYKo/WWrJ9utGdzctPThA7BC3el2yCxUrSWDCHTxuOddbovSn
eOBnCjwidTJZAyNqvL3UWUQUY0SVqyv/KNIwbVKOCzDMKo3bs16Twtq9cCwfgm/6
Tetw1yCEGPpXSXRliGR8HmjYpFrOTq0GAAywcn73RP5AoEN112LK1i6vmqXksDa+
IiF/wfmno7BS+0Nc9n9RwsYXkXQFblwlPpG9KaFBDmkF7YiOGxQm9FZywKSFVfT1
bWl3wRovJV1pTWp70qnbuA4zMg7x5NhvfAa5jxyrC3Zq4uirO1GsD9G2c64sthgY
dFwTlhqCsZuNRexD+GUHLm4En5nZv0EcA2RpCBSbz3j90+PJpHhfmPTW4turaG3V
3z0OBmgIh2KwPfzv+s3/yJo+S8uQx1ZEqbAKFEtmwHD2vUFAO/rOJbIAC9rGi6BB
HP/0tDt4v2QG5xv80mhG4Iy0jPFQlPB04TquST2bQ6+sDxQ3wj4sykbAlEoPFLgA
0nG/iG9mjpxLaGxJmoXF0q79Z8M3VFs1zRXeglXSHxPSgcopTaDJJK0HkpzC9OSO
s7jbdWyzDA1hYTTi1x9DBe1FO8ZG5e4JiPvTEpHR+mhVBYEBpwZDtCenmtyo4vqe
ljE7sTLP2nFtrCh07P3KUfWZkEW5P18FEYhwoOehnjKTEfAwpHsxtZYCyLZFMMj8
5l2bOAbdUQWlGjqSAT9lsS55WmYh2KCEWpa+VxAdV2OKRr+ERtTmL8Ek8Anp9B0h
k52d5d1txHfZ6aW8DuDsl5iV9XaC3ax8Xj1HmMUHe80lV4IxSKzJ72N6bdji0fUE
Fi29zPI4EiOjV8q1VG03SwTEzak/INJKjPCGD0W49aPMfQoDFaHcnHkd3TruJFvC
e+zB/QdGTNVSqlrguORZSWPC+Dr0IWz7e1R2peSFkabR5HIiJRWx3gVt73ohdb3m
o4n/nRYH9MGFZlCOhltMco+zoW/hXEBPS9cXtUg9Zr5q8ItVebOrlhVoG0cR+FUU
6vJn+lIjPA7LGI8SvpYqsi/INJP6Alpu7Ksnnf3tV1WpRURORmEjm6TMG+a8kVRy
EgdD109nEh7I47BfMx09od9k55Jo8rAW6f0ZCW8Mg491P8QuSq92RQedeCe/9gFM
Ev2Hn43WDd1+gKJ2dJzxf5uRTMGcAVoOGEhAd8idO1WPNaK0EY+EZK1qoIZ+hirp
2vDQqDvjqJ+D7MOD/F5rN1bRcOQeB6GjNmg/uhHyiv1ziV4gzBLqvvgBRmySztrM
3Jeh1wiyyfFZZbcH3W8QGNikGujkmzPnBPD2EMa8ruOHpcvCKO8ni+vL80chiXNw
O7pI2hCALVcf6wvtRNVSXpovWhUnU9C0pAuEikJ7JuCEV9DfoHPcjAq/gHRdy5bc
0Scvyn/76jBs+vThwxSqGXdKPdVdyIC0cezw6HKJ761l9Xq24Jnf7W6HkffX+O30
Kbb8Rn/SS6nyOdxMdGZcADHdBVQ1DgS/Z33KwdYFjksJjYFD1wK0r004Di0J5AKp
uvdlOhjyV/KjA7JJ79BEm/cnCn0i4aEtrR99MTYns/ecYOjs3Xww5/aypZ8GQ7W3
MkKhW+ZXizjpIWHFI9vdD+f9DztLAlCp4d/Me53mnKbhksMGK0mQbE+Yy9P7Nx5Y
b9wiguJekR9kub79fOBL+XH0kOtfiAty4zioJFrZsoOVMmnmFJL9qrbE0RAMA+r8
8m8k05I9BypThefKc7OhK5IJuHZW78vNRAXiRX9CrkZ2NXk1JuM5gLcJ4WtoU6cT
2bl25G9RPOj6LXLCD0Gtyu/KbkHvR95cDtRrrrFxZYIC4kzynRLhtK9VNDBvfOkP
me3t8Bzaa4/vlaJzdxuryFwkfNzDSyhp20jxaOG2VFqzbfuB3tBQ2U/gj+6pl4yg
GvxI7UvM/CBnkigwPijt6b20/iHBzOOsCjZ8qpVw5ON36jdJBO5+0J/olsPC1HJ+
akoj/X41PGmT94h/TTgyVXfVcm+1da1/c5VvM4CF+zKOIzuBIc8+ZSnnwBtwggMX
I7SgePPFBwMVuxcpjXYROXL+l9HT9iLaxhNLa7nJTcNw//Fydj9UTNdrKDQgW1Sk
+ZhxjKikRmapwnDn6efWT6o8iEXJ8gaXDmac1sLtJh8phhvEU81GbhjFIrUaYIoy
qKnoljp1P7a5YiLx3TgMW0Lqdy6sKcABb36nemyFh/YDO7hNX3B4J1n8yQlsuaaO
Esxhbie924Uv18heamhgoW8gdedGc43VDRKeSpHpArJZbGQmbZ0zowwDWofw3zsY
l8THyEkidqK9jVCf69OKizu1JEkdQrFRvhAwmawbHtpv/inq2s25G7CrUv7g/XYc
rrPiV+IVBTZv1xFE+I779hGRdAebV022hbg3//dt4dTkippVlv9961pc6axROg9T
k0KoT6kufIFbNly/tcxyiqsnurhs6JERotafa/yfcBec2F6gdw4njVUeVHJ86V1u
W2VFHxYxzPyKOMslsRfLwqKw1jneJfB5WD2UcIEfi9NaUGcUGYVX0cy3wv9FQu8A
nkbfcd3zaXe+8Y8FNMG3DY9NyIH2/n/fjHd8NfYdYGP3YgjqFcR18sHktNm06e+O
5+niDtylpq2Z7XuiMHTdPSpaomSq/jsH2XOnilvMNHWoyV8300Ge2RjB1zMe2EgC
JH51AUYuWIS4uukE4Np/B7QUVYruw4z4qxr5T6wI8oBqvLn/E6d5uFqk1UfmYm1j
wAn/LbQTDa7vSohG6iX9FcCpjuaN8xkY+12YMgLTvtAs5aH3j/Tz0CGgeZtgVDSB
o2aaC+UF7MRlH2Z1MnwgpYCiVBCM4A8rSIfTP2rvO011G4i2F8IXSw7CtoEH7Npo
6IEHJNxJLdCSnzexJbRhcdeoouR7VD+2y8qBqe5q6i29hq0Q2qQD3c8TOEWVdZdY
W5uwXRHBQ90UN0bMuS2SKK6zBrzVxC/ONyDiRQvcX8fpJr1WLvwQWq3wCBHn96Yj
vkzGgXkHBKs1QsDf+iBBuYLvIJktXzlL4o5EQ2v3Hzplg0vU80NyQzKhtAvT/iCi
/hyFgfI21VKqMjQx9cDfLJ03RtP7zFmPV+TarvEOvFGmsbzrjXV+j/QaBhaCDnkW
yvdfsSSiIuUPEt2J0fZISRrnJM6ElhTInuhmwYsr8ZB7ZbMEFyhFJdGZTdUkJmOy
vfB0qwMzF0kZki1hMzVVJ7u2Z60FA8p+RX8s3m1a+/aEdMFNR72bSELcHdocd0D9
M5fvLaXU9+P+3cjAJyRmjqoh0g2UIMt+l9htE0f/Tu/IuS3n52SJHvtwV3z6iStF
+UDSYw6QW9QHTy4b6HCqghBMKkeKdmtp8m6K5/ggJcqBooFrAWAXpdmsVbm2KdXM
l1BpHA5O1nXoOFgjeLUz0TStC0+SW5JskFo2UcOH2on98THLeoYscEmblHugwuHp
W7vgXlrtVczmLkfsY7HPOBpxnAY1zyFFd5dLF5sz0LTO0/jdwVy6bPsL+9O9nmch
ZMmiUM9ZkKoT52DshH4XCORgQIoQmEKVNpJuLeRHnX2yhY2JCzDHNASlQDACPwp2
rvfFyqw56iJOr480INfXgpS+WtlAQIOcIiagKoUhDSmlaQdIra44jrFgdPGRwJbS
3uvyt7BgvmEYyGwzDFFmBLhAnFoWD+ZACLgIzyX5mxOrM2zROApzlNIlGSMULos7
Tyb+mHwyq2bKU3AP3Dm7kk0t2QdX1NGB4Zf8SrSf4ht8+VqASj+ItmAjsUb2Pgyx
fIw9yiUBwFR2PlHfq3kGLGPYkJ5JWeUF4RAoKCZhpCEX/W/AUb7DENmtTuANelUU
87PU1QNkQCnByEjATWHhGrQHvh+tXqnoG+ivh1Xn7vaPL6b70uPOVPh++2r/KCXf
ayWfkSqb5RosEvCQ7+8NRAbzykCPU0PlhxjPSyI+2F08i9+YHx//OXSjvGUX3e2t
+bFCS/txZm6eGwuzY/7nDpRqMsk5X5U4uES+PBbrOjdovQQcy8F8k8HTtYtN8LAi
SulXSehqC577pb/dI5U3wH7ddF+FlB1xPfEKavYeR27b2LI3mHaYZY0RxxSwcXbD
99COf4j07tYaWlQcEvmV+G2+4e62BJYTKsrGuF/vGecSJaO8VBwknxUzZyWLtJPv
MepcR9Tx41T8BKD38TRen0PYEe3iZfSFBiYXTuwMmK/mIug4pvifYkp5lMBSCjam
7KnDcyhG84z5IDtYexnxR/AjHpDxUlEZuJ6z8Z0jwM1i95O8eJ/vtmM8H0mjOH0K
CDbapX1itn/CSQ3RT9f8bv+O2sFFt09MsfDUfYa5kUxki6yNqNUf1J3wQnWiHdBG
1A8a/hh+PzfN533qaanS5q78seXT4CATEbbZeQlKlxTezdlL9EI3BCvcCILXIp1T
uUpqGqvRZUpvuZEa34xZpYPykmZc59ssPCtgqoBJxYYqlM2WWgEP1rzs4ZFJkR6P
TBX55eDL0R91fm6AsB3lfUByNg3xSurcmQ9Z2FnL7mni0UB0wE8qAInTSLQAxGUw
YUifE+EfG9GmpHHPHvXACAxTc4YPssTCJ6SwTL2eSofqsuMYkmgh6MRrFWOzQgeB
DTDsnxV0F+JWMEFTeajUOf6Dk7pYoM5uAFSXeLn1kq7sOAOLx/vDvqEhLfqIse+K
/9dA40kAihrR7BKzSdkhevxfbGyu8vsZqm9CJSYvvVJ/uiw2nKwD0TvLu6BlVHc3
IkQh6oZYrpMvqaVI2+CIEpTn0hFvYj/jS7vo3oWPAUS/rpY7x+p3I7T5T3Cc3/an
yD/CgYf/bNVBjakejBkvXVz7QEIG3Mh0SZ40y3QeMPWm7Yc2HX1I5eWXUzHgEj0A
kgBIQ171oZEDkM/ZRzc9l5wkO/MPypbhv0PjDfe4KgYlwtdW/8hzlR0bMj50U8BC
7U4nBiJSSLrPCSVwAp/noIVUmmGBhVfPSIfF8WGQx2ML9ldfqUXma2RgpogsMapL
/Od74yhnMZ5HBg062TdfTM8avZcIrjJhf2mOl1egAAwbGkB2DCzbxExp1XQ8CQtm
Z2u9aP0Wlxd+aD9oNsxeumxIHH6QJTdaY1emfVOsV0ed2B7nq/nhcXL/aoCby6JB
GXamQccXRcw0H86AxPAm5gOevqY6z0HB7bGhwC06UIWtqn1vHElXP/HJPH/Ccfv2
KgvAmN/beX/T22FUBuxv4F+R6TyiQDpOpWe2u5Jeu6m7WkA9j6BynkfLDjGJxG22
K5Fqc3bi5STkphn3EXYS9GO2WBaoX/QTkHidYOV87CQ3iQkGh81lM7/O1rK8J57M
4JN0AZrOVN6jHo1fq0XKZV2sglgBqvgbWKLd5JO3LGLiOGL8p0Ic4lz6vQVRsK37
a0ctEur5RfjTXIuOIaIpMW1kenBpN/rBHlxv0nIVaccfuS7XB6ebJF3R3+ZGbuJv
truR/IBSicLxEc1IqwD/jL+E49WHRqr/508uXwD9nHIZ1H4+aakNJ9qNHOjb0Zm6
IlLglAco0awehibNVRDMc9OJcrqjm7mRgAo8X8jkIxysVoBp2Dnz7kPl2Sg3mron
89/m0W4kAe4ad9/BsuJKqwBSZtmxO0eoHudBrhZ6CBhQWamuL5vun3T5URBdLT7T
NrMA4rCkGDx2h1T5W02PtAjSOnrMFi63d9VB4G4EwFCU1tpGRkgqSnGua+kgwPUP
6elS1JU7YvMWQRpyqyiKQYdrohL4T8hJXq1lPgpOGG88r+75XM9D6wFmhmdt+H0S
AX1bMwtGc5yC+ZHqcJEzVeJXSqFpn3LeWTTwCjQ1m/BjWB1WCDtPw/0nZVoOre8i
0VxILVFPBfqdnVH5RCxz0nop4u0SARL9LHuuaj4opmjNQcpbXaKC0ljmNn0f2NjM
lzbwdyCbGBSHdjdkZeQ8eZyH9heH4wo/tf6iO02cEAZ3p+JEgcWat/2U+0vwzLme
iIFRIwreem57mQcEl2Q86fU6Bcc0+YsTsiZyOxHrNWrVhRzcnjnDUYPY8aa3MdAC
nEJ4KjxMzACwQSn2fRIzvSLThz40PMihh5jj2luxzxwK6Rf2t0hluYEiXsaEuKmz
btZXWfwDFzCwPGoW0Al4y1rgpn6Y/AnAD+A1baDzFKl4YI/MW/l5ec2LGdoXvM64
AZthrX7iirTVCD9EvXM2i6m//f72ubhdH2X52P9jLONUdPfbeY1cn3IHKlhWvisB
qw8cSaUx6aZ97uUKe2p4Tn5Ijm+vAJcP2m5AHpR2jw+e5R4mjF7SpgqPDjFKnkN3
Ralz3QEDNNfRjp6885RJt91S1nShiRPdx2v5C7NpN5yP1f3uRZgeEXWOfRqShCco
ICjn4C6OTrUSEOmUqYt+YPQfyvxA4ovFBkOtI3neIlVAxClnCp7E1rGBSn5uQCxF
AC2zkkzobPLBEtWSOU4IYeKxBZR+uPYv5+1uzzcHGY8SFqwvXVCBsMzQGMW952uV
PbJldmkcETbHdEAXadhLVrZXjqwduu3239Vc2VNXO2gHmKzUw2xMtxcZhGaRZZ2M
14PvRdDFeOwJCKps7Utvypzsu4g4Bg4QsvAjbcH5OgvwqokwBPAWcucJt/FpwRIt
E6FWMpYJRLu4P/Mdn7WIoCuHGKuoTjsh28zz8VoX9D+6LykKKlXgz9RqKd+H8UI8
3LetUNqr1CPflraCzxCKU15KWd0nMHqjdIanBXpqDv0a5Wg0xsWCc4n/Oxbn16+Z
PKbj+PRAgshBHPqSO6csmUZus1eHgiZzZzZ9RA5TVxFhfDFXdHZk6eaNcj7YVO6b
HjR6bd1z+kOd9OXqFxVfDs3OiZladd3rf57n7T9MdwuvMb4ghjV5BFDMBYStIUDf
AXImY3S3rEB572y8etjn4JFK6DOJL8rBB6Jr5ePGcsC7JF3A2Ol30rAMRWqw3aiH
TANEE56tFR8Bg04JsFHw+C6oq3yxCht5BF2UTuQzr0JrO3Ec/pDdnrk1S473bsLZ
iQkJuToFbyT47XgfYucmtxnGX8BT2khO7itMdTXEy4iiX/+VFW+icgzhMktOCGzP
NfqMPVMtUnJ6BAVqwzWxOWzZ/+hKIFbbxOQgWEXWlwEJkqymIr6p9D+UB9uPCFi7
t6z+QgAitYiVQBwzFFm386yzcNbZnX0ea+q7Kwine0N+IuDzbPLEybs81sYbcSwV
pXkmneSqaGQR2B/1ODawjESMjG6kWf6hcqRqJbXqgTZMQaheaSSoguu600Z2iJ9J
8Te6xsoicc4oU93VuY7dwdAeT67VnhnMsBqh/GcvDkQhoRlmUVrTqxiDAczcrtc8
aLpoYkRJ68o98QX7jkYOaWDXwrl/kLj/aDouSfLFV/N/2X9JMmrv4RacQB3BtEGR
13a99q/8xpye9Ml50bbDIfjOAmSKjeIVYoHnpQ6KrO+vPJXF7HEz1BirWct9dWt+
tWnqWFC1sHuqTcXGxIBsBHDUwT4z2r28qOTYVeRgEMfAs5KWPf3+4hG7g0Gd8yMM
BsU+aYLCJf/CBEHOMPvWTY4a9xIs2H1Un/e9Furrov0vVP/9XlJLeBzjb4RRdbs8
bVFl4vKajYaDlSNEykZ3+s4cJEiOJIJUrwN5abDTlFMc6S5JuXbJKriD2pcPKw++
SJTbVcoaHPf2Ntb3rcD8U25/kL64fvezFa09tVVYjaK1/DvJfeGeajTtNYs56gUc
YAPm0VNO6mQr0DBuCG470UkbKXi6l3tUnz2+4fTdHbFXIlW8K948TIpNV2ZuZnYg
8So1+6nLsmkk8D7+qD8PXpkSVaWjyTMRTVGhVT85wLElYzLjBmdOv0CFrhMyoouZ
XYLunsuXyI5tNI7/tQsmMyzg37N2A6m8hdDCF0cr/Bbhd5CQ8aLBZiGCIfkL8eWr
58BCVNYanwC8tVLgC0Ey64SlmsirN4K4DCUwi8l7HUQ1C0JELhwR/36GqZppLTdJ
Zm4e32QaxszC2VLqFEkp/M1sbyvBRfimdypqfmATwIxqRxJ3H2EuCqZvUyU6RfCO
oigKOQ+cQrY0lgGUXANciYlhl37txA1+E6uEeieWqk5mLMzOUOjxydC6TEmj/A9+
550xG32oN1hLlMs4OswWTxxPiHxgbKEke4q7FrBiM5Ab1RyyjuCy7L/JesgGrxY4
dzPTi7Z9m4V88asdJeBrdoUlJPRdayg/muuBI9GsXMRC2LEIHRiAPfzznU1qT3Jw
kmICOpulvt+kg/EIu+9beJc4cPrhKmPrqsw58UV15w5ZE7iowG5QUu7dOsTXnljv
E+mNqr9jnq5HGHGLEPS2Gsz3+qyUCG2RaIEvZefIm6UViUbCnhaWFwz3yeusAVN7
UuOF70GC/bQyNRVJeMqk9DfywNgWfC+IQb/PI58wMUlERD4KbRuak1CaNiKt4Tq3
mUSKlWM4bvV8dyVlnUytrsJlEqrUae1wx9uDHVerZgPbm5OA8s/W0LVS5YEYG/sb
oqHzYb4P0CQtFst6lPk94tQ/8qRHN7QdDI7N/gLRfUFS5fhpM78IiEepBtUD++OD
HRzuWp9UU2VyMfskAhTZZFWJX1/7WF9hDdkIb+bq4uQ7NOGILhEy6JPfoGxq+SS4
cvFlQNInYWSSTMxW5a59AxEG3FUFECV8aKjPzJ+b8fP62lvJg5OQdrU8RAwYckCw
9uPLouZ/NlxT4SBqAjX835A3bPAnscaLpLOysxMVXJA+JBkMKgBIrvK/aoysIoim
v6tzEcjXCViCXf165DqTWADhVtSV2pylup2PX0LT9P/oOva6u7s/rVPTLQmFc/zw
15I0w41X60BCiUw+9A7ZZREsFSz4JZGG4DharhMJwGJXa5x3qEPyG3OfCU/eFHZ4
UxeeFBOSNDKcl/1rw0IFFRidal7u/Dosoq8TlkpnKr05im5U0LrN9/nFo0O0+QMa
+8gLdXAQMAYQGjuBQC8YRYNJx2a+U9Tcj+VXDFepzlZ9ae1pYBy1hm5Xvj1xDgwg
eDvH1tQY36wnfsdLqQXCVlmAwB4uLlsnZXG7+RMz39rk2iVb4NexpFc6WBWJ8UoO
g33jiZubta4pNyqNG5qKQv9sKsAe79Xq5X31pKmbBqFoxI7rudkWa2SCCUr9Rpje
N9lyZ2B6Hk78OWfRy4/Rv/kjQ9FBqumc2Mj52wWqCop0xwipJ/EvMydpb2ZZWWdF
H4c19Pmk/qMfuZMP5m5wXMsS9xdKgAoPnzORVVfze5YOd+C97Psf6JF+SzC+dO0r
yqb/Sx0CAv+s2oOnF54md5sfTd4jdKb4Tr/Q0Th5y3qj0QyOH8JlTVEJGQu4Z1nB
W3Hl8HTS78vDotuNSbWvzTtr7OxJ0yKwq1qqOTf/oDrHxRt48jJQnUleJr+VdDx6
jLpEUyCAcVMP5Rq24tjdAUn7wJ9IOmWGanczJXAMtnkMGQdRnZUe6mVGeoL5Oz/8
DgqaQuQup0ODxE/Zl38c1scoTfthHglSlqMo3L9d5MsKn8eGFvinXlfBMQJsJzNg
hmAyl+qsy0T/NV/ZqyiSOkb8LYmlz8oWwP9t0PU1Wnqp+2DNIVyx1njCrGG1qZgf
P3PG7FVt2cIGvsNBJu7xH5DE1uDMwhHFTT/Zi0F9CHA4yPhReurIGUWTvzVIZbVU
L+nPhJ2iYy6GolkvtcwzScCWnS8hFVY9oZTGZsYdLDo/wKQ/33NC2TomsbQy6Q8F
YQovuXG9LRbBt8ZufSmZ8ET72YoAFfT9c8VunjOGEGHf1v+PeoeX4XoZ1HAYPrCc
kqr1tKHCf0Mo+kPnEzJkRt5xlfDAtCHnw42nYEX/mwtD75Lg2gz/TaGWDMHlrnmv
jHrnT5xchdPcIayN8gXfoZZujCETsZTHCPVHq5niYSUIa7yPjwwN5OM3zq0/LyWf
ZiJdOtpy0CFxS5hOs9eSZ9EZM2VUYpjs3kvpFR8/pSpdeP07/9LWHHxitLNYIp/G
+nO4uQabzoQAHhDkN5GUKi8yKrsGS5xEvnWf7LSLnSjOwe0xKeBOLvllaTRBTye9
ytvzynBj+mXMCvbKnlUWqTqpBrtjGW0RJ4N/TEkrJVITFyr8m6kiIg5ThRgvv2hc
z8PVAp0kfZtq9+WaNZfVb9+XbwLio/rjHB23gIIDq+q6VWsHqtTVizAM3deWRtpM
E9MgxKVAakMSqq3WGluKYbKHJibQjss0gbtQepL1Q9YEqxr98wxCwzMkDKdXcYJE
CTgNu3YEvgRXQoTtdsSoSvXkhhyT0XoU/YppC/g5n23QdVpADazpQK033U8ZSFU4
lvsdRb9G52nHXCDDzlmvYMVx+1qZyjnUH/BbJg3Uq+bCbfEI0gKbwLXfQ+HePuwz
hSxtNOEk+WUSC319mX9rVmKOnEdT2bPdQbKZH5yx8KD1OuHZitNLYVohmELNjdFC
m+LApjBtt8H7ZLtMKhnzgVclGG5keDMrLk7aujFLSqsokppYrC/ekiATaWbxY3/Y
5P+gy3ZhIv8RT5m4G1qlE+cEMWWwNZNOQ/wyf5B36izUPCpK5Al0DhqoK/DgsG+M
xAENcb6IHq+E/Qpa8M3SWzt3QdKAv74yE4XOJqosCSGmmo9ucF+dxhNbLTpsv6q+
bz9tKkLCqRw3KLCIU2kNQn6UJI2GomBTgo97Fbep1npUTTRFIWzUbVArlCB13Pir
KgxB7AhCxg0EZ29/qPkBUdnEgyircDVOY6wCunrGYYPisoCLsYVVqySxxDRBKCs3
lK3Wl17SRSX8fATP5m0JW/tYD81RGN9zS/9ysKkdK/298vH3ul9Otrj8ugaeZMC2
HlZYvCy5dC2IDxt6uFW3P9ZVVRM6oz4OkU3jcSgWWKJl+qu+bgt7LSPXKzwVeH+E
9JhE2A5L7FtWpqCyZIfTgKOt4TOOPs6HmcPAKItKvuenuk0XhZ1r93ZZXjgJuU0b
HT4BqkaoMdxL5uxfWFDNrpqUp/uYbLA5OH7Pgtn0l5d9ibvXqUCkaHG6YhUjHt/A
vnj3s4j079MCSFHAqeCEqI61tbm4OiVYvVQdgMbEqn4YTOtGydH8eNiQsJJjJ6CF
TC7vLYHMXBgD4VMVeF1PpY6s0vlZVfWdGappqLi0YfSA7gYFzObHttd7xqB4KRjc
6bI+L6qgqnVrB14EovrSP9PEhHSfMK7LKeOvgwOT3rg2LWNC0Ae/0EjXNR00yxYx
dPweP4sKW6vs80oveBQQgLDf7/4O4gnW1zCkdHLnEcxdOphs14gvX8VtBDl8ooQm
4GGnlKNSo04nZuMFaYWa20bl7PEsrNOw8yXOeJtyWEzhJm4q/o+V4vg6SVE3mvIe
7s2LFs1oEIbNIkxj6y1QLu+PK/YVL+CCmOnwhvzSaXs7gveZdm81wtVLORB29nWT
/4Zq2hqjaQt5NTXJFCulPr6OLpL7cX8bMvHARRg+3Nn1cP30lwvACQb+jA/Rubnu
LhtDEuhCcKgQMJaAhyeqI9U8Ap+mfuPCOkQJvMDgP22cJFXNV0Y5KWR/fqCw6ooh
D1HqF8MZrlV9uA4vkMKc8Hy2GskRQMjtBX0PgS2RS+atu+Rn5uJHbzDs4wN07IMb
rPQhIL67Eo/LeWdlOokeE492f0O2EtsNpS7g7IbmpqYKZXCKIGKGK0/1//pAV2Jk
oHFCyOLr2CrWAI6Fd5T4cgQ+4cv9C7OcELJY+kvBnLKOpxymVhAE/1dO8EedLVlU
ZdrmPt1t0MChPqCae5752KNkQUq83UikMg9n4LXLD8ZBWUwc887P12BzCvFR++/N
y0AfovFm/KpMfZ+4U8e5HL4pwI5Ph8cIXk1imxjQ/Nuo7r1cU4Z37kA4x97faKQO
9/v4V8FzDDmZEF/FQnIr+5Ma+4L1ONpQ5oxZJ9CZ8KITY5WgZ1aHWD9+rmb0rdV+
ETNBZC9qi4ehXuJDj39ulgicnSTFTB5bKoEefCYGGPWFuO66pRVy3rW4DxYA2TwW
R8rrfhM3yfIlWhAj+KVBsWy06yfAvqUAWlA/Kumer3z7CvxcDUd2WQgCOyV4jPU8
jDsILORm1R+vmAtbBo7jhrw+r0kJeahgFOdkyTa7RauKNvavytPpFF37Cr6/6PXo
w9/jwoewbnDJITDgRwFEBNYFHYXJWtnbPTxvZajM7ucAczekS/oKN2MFkFwkICJL
PKVubNxL0XEx05IwphQ29qsONiPXOlV/SRvwaohCiFjv9a/J2KF6UxRViprJybu8
DLOHllT7f3HHAywz1joPfb/EOE9D1sz3I2wljM7iRdM0nE7s9GSZu/ewX24VYoN8
GHRRvaio0R4kGtGEQQDKFpYbi5P+2IFChvKamzzzviCLXZzj2xUy/dsyQ3PjwugR
HUUCgsr5mDKcLYmqD2RBP4lyFUuhei3hvZzJbSIz4hmmt31RhqEIiqd1wa0dt+w+
w04jIpoZoJllS7EuLwWQZRg8XpdwB/DnPMvVIp0yvgEsqcZh533YVU7t/JryWBh2
cG7bo99qf4Ot+LLYZFHMt6NY01VEIfh1qOzkCXxsWy/hUFeJvsOmlRRzVZnAkCyp
5/SaRiUhr6eYM4YiZsNQ14cMxa68bwMCVgurwM2S2n7b7S6HBqVMHQEsLijp9T1h
S0no5HhBqf1n5tgtlolg837o4UT4JEe3TyQgXV6K4lnC1zUwaG6jzmLsyO9HM0th
su9mUMHFmq3wM30v59pIQBMe/soGZHXEs1aOwPkteL2d/jYn5kzFq6x3cvD2j3aK
3IzIXJbCRELNmO6hfKDQsZ8ufWu3EtROxLaFexA3AhUMA61pzU+ImHiTBrx2d6Ey
VtmDwFiUpaRKQ9TPLrEUBbKPnP2/an+evJoDROuHpQaqSxsBNhrpA4ZX0p2hFFWt
ckDL7puJRIrj8rQGJM5yzfYiH54aBVcxXbVmYpmhedSQF+fdytBwY4iHDwxdqpNB
/AwwxXJjHsVLLQ2OYykWxFt0ezmtvZ5uF8w9e2eQ1Jj0Nc5L4PWicjFzkSDTL9CT
d42OKtwDFs4hwpDw/FM5CiPZdf3/fEQRYVeZqnq0OxcU1S9sxRSwBE3ULoqE0wa0
1DyLciUmFk/aTA+XcoFYBAhcbUusm6g/QrhiM9yzTleJYB7PCgJ72FRxa3CxgTIj
EfxWlLidVE8AzUgfvL+w+8hAddY6dxQHul4ZL9EkB07dvcQGQu0iasZLfCzXP3LM
kzPidYfJU0eNK5kV+QTHMZuzKUBk7iMXMrc8RGAXE4Hc2CDL12FS9HAPOMXXle8B
qh3Qw7s/rC/8sgy78bjAYSqsFkY4E6OQatZtV02Er0tdRLYlNfbRwrQORQQh3jpZ
aOUvw5vED9JUtUG8G3Z4nc9WGafZE+QKoHULH911uc2IKI9kXuE2d/aZwVdhxl97
czDIgcsJd3hAKIL91+et3Jzbqd0pF+gYzm2qS7vazADZNMTxXvNVZvr5N4MNOKJl
PIdyebbh8VLwX8f47rPKkda51Z0SOqWyY+VBWVWNa0xPeMEuvIDBuVT/4W6gXEtc
7xh61nXRf1uTcF3A8TmbYV4aoRtevWQmLyO0azg+fWRBvXhhhKa9WuKuWfbKvWaQ
mCSDFpTZ3DBZYQbIpKdUYKNtzS4gfFvJ26dSKYq6wAKFa7qp/1340HnkUKLw5Q8c
T98pggKDFkFUtBmjUyW5XqwHcsg4j8fR1S0u/tTVx5D04I7MR9Uwe2zqyy/7JOLS
/ErrSUtB46kLLLoaDMaGi9Jb0azdeBJxfkM7Fg7T0n2yECk4izwA3AKWw9tO3ljM
MTtVtshflMdxm1TA8lz0bHAbQ3S+FQhMWY7Wt4sv0UEALhA4mnlApdXsGdpD7GcN
1iOzgzdg89X/JXOD/xImU5DDhQRtbZefeuizbqlzIByjMAAYCGEHBucC4YBwXzIv
vLOSd5g7/1rVTHHVpf5SGmyv1U9hpaOlCmQKS81uS9tgPovGV/K0InqgxXwglRzd
LQqDJ2BzlTgXWdOtH2wwIeulVXL6L1IQ7OgOSB5387lprNJPzUaNMnOPUOX7p1t8
4h1b06inQTiF+GmhuOrC7QSaM7ghYoVtie2VSK2UrJgfDKf7eRnqTi6SHmH1AZ6c
p0wP6T4aHs3zGGe6ImSmDAnOtBrtQSm+zqjurzaSqT1BzfxOh1SxEPybjbkVJMBG
QTUO+m14YLHDClV2f+S8ShFMmqtl/olP4YqwWFsz3LbPGDT30s18MKfhsv4/qlLi
DBEMobejpBa1ETWbD+2El9rAMMLqDSot2W7Z3myumsfW0vKR7ptyGd47uHWM+ESR
raEOmSx9kY0TwK1NEnYjHHJxPeQZh3Wp/WhISvdYdVVjxBvkZ4JkLij0SJSiSbKM
YpLDZLVhiUXhPuNSu3V5h/lzQwmC74YaYWEZEw+fucF3AxVLAjRP5QoSLFHWnL27
mwx9fCXNX76gZq01ZzlE9lDeASaIRLP7A9DuGEpGoU4wZEWpWKDDTT8i5GMgOqoT
S4+q533q5lxjWBF+Q69y/QpDoO+5uAQnmFF7LYmWSQWBJOMDD6Dc5F4t1z0OQRsh
zqBtiG5VVk9smiEhJ81lZqxxXMaqDO9I05bwR899VSZ1Yb+O3k9WILKXfMjyqg4N
RgrVtwZ1EOjR5lcm+WHtT2j7hwV39tmwbWOGzVtF9ly+dvBc+alTAbNSxAPL9N1O
g4iu7srroCsOU6Xc61oWZQIR0l4NiVY3YKC02FXB3pBMm2DNt3rgmCnE3K2WUDbl
CfY5TTqQEQhPx+sFoQIf7sBegCjZGotCVku2LGEKDArQkQMA4RwgC8+PHbPhmCXS
DCj8xIf8KtsJg2fSITjknoX08x/hjh+FmsZgfcFyFpdoDAAbNBrB4AZE6yMGLU1s
lUjGDXw47q8dHRgKwF2BJLqBF0f4xMVsO3c80NSNRVDbVUTCVSUtt2uzdBabYE3L
hIX2tlPs+GEXxq759fUyV9kNOmrtyjIxj4nBSfJLGc/dUjKhzJw9ZMCPHzjqMgkd
DqVkl20rCXjYHpk6HXXA3WhxR+i8mWz39fknha/0Gl1QO1s9NTPuD+i83qfFmk21
ICeb1432NEtUy/tsWVdSrxeoOCKjssJnp+MeSUtTb4uQwE2TpegFE70pd99jUM6h
MTk7O2rjCuEor9PMPxzwCjuSu6/wI91TZ5/xGgjsZzXdGIHzDk+UIslhHVUCTHtL
8EzDb3PKVNSJdUbYxSYnvE8wg9CZxAClAtxX75zi/AEEYLkFu0mld/3ktzeOcoUI
jVTGQgAOhjTTKsxA7vmq7wjvi6442WeoYuIjCjGCA3A3CErkV82zymxFRS5YgvlI
rXCHET1KX4sOKUmCXXkSeEw15PJTPlUxo5LXr1X9DhdnFzmeLRfyL8H8rXkiV79J
DMTVuoz0/60K1iKmry+ZPD8wLtRC/xU/kXAiEckdGPrWov3Ovz+Yn/NRi5+Td0Jd
sbthhYbHqotST5zTt0h+DgyModtQgDZ61X+1qajCr3nYI0FIh6cV/CMBTCtNzkur
mQii0W5KGtAIXeLclYvLtrue1loEU8S/cpq5JaYtxETkSz+MCBiNlbwj+UJVU6yh
RXfVVhOsAFIS1URpO6kNQ5V0KC9lTd1t3vr5AUKYAvbG5NP1E+Slk2mgqN0to5r9
vu0xlE9Iq9zUxrP/1qC0NozVKd/2zleTkDlEX0nVZU2nkN3VqZ58VlswWwYErKGw
eSyqC/pB7UiMP8CAL2YW5r/DYg4nUpfx9TeEfLquWp1w3fhi9h1/X6ctJi5iCx3A
0tbmED2AUBBDrgw5Vh5VvMNvgXESGuazHMcSBOofctaF+KEXJfD3kKX0YQ8DTdmY
m4VccB5C91RWw8FYiHUEyv2T3z4+CeSP0ppDVCOe4fsY7kc9Rms8uOUoWiVlaur+
zAKLP8KPCwoiPF6ZmkG+7mxqnr3uwfNm1m7/PmBr2EX/yflD3Ej9sE83Sd0H30c6
t5SHRzKu4xtZY80QO74QkwjFO9NqMG10BP9ELu89u7v7DGSzlOTA0l7BFX1CQPiw
lrtPN4AebkFYEhDoQcKtCa6gTcwCL+DBtkr2wjJkEW548cSq1XhXn3nZfhult5e8
IPR3vklnFgruogGIRPw1WcEXTbCVZSiNoZ4OkBlH117z1pIz3jTPb5b0e0Se9Kx0
LBD5fdLerWHRflzVea8Fw3Kxt17R30gcFs/Ze+4kXhkn0Yf7o41hnrzRIBu9jdnS
1iP4P7Kn3LD+Ozeu91sDiG/lXCa3C44g5p5ZsFMtDA5ayVVKZC9B0zQK/+b/9PYq
/qU2ADbJtgj7ZJLBJJKqW9wk7qQZkuQLIvGSFBBqzfzPVOpGk+r6CABbOA+IY8ci
8KQ0CV24yWBk6Sg/mrswkOPj/ckFdjuQETRPjeOxvwmwW+lR6u5UwhxwtKivySLf
Ljzw07BxBzk9mwpEfoOA4lJleVvOTBSXGLzIGvjDgRAbS7zGMQTVWCNE4nJpiSm2
GG22CibFwjpz2jVT4CbcbJB6JIOpU/bDpBXZ1N083Jj0wnUnXb1hXJilCYd0w3V9
IFYPEeAffJNaJqIUj+oz63pPmA8btF/PyRDzn4FnT9Gm/XsjIQXOhT6X68IvlI14
hJylLLn9spyKxiP4Z1VeljwxX9pWavtDfZwH2z71EYDQDD/OetnE1C4Z0F87UGT1
f8fK2e3V3V8uJOIFme7GVJt9oCEh2gPqkYUvnfyCpQ2Ll413Vj7n8o+PPTfHEeKN
xNeMeib8JR4jaZkJAuMk9X62utwvZ27jSEhS//sKlhmJBWJp1dBooi55xZq7UP1K
c2bU1kwz+omo05h6jdqAeadHgsU2RixxD/wYWjRDeKJCyCdJAB3BDlZCUonMUaFG
nawKUeeZZlqsZ7UEEPpJ2UkRdWpemK6PgwBNxYI9FX5ouSFC31jPXOdxneN0L678
O7YToNmPdxFQTHn9LU0kBElBAPR6R2RvgMNBBKtC9A94Tk/IUVa5iZk1khWS3X/D
fjXj/KpWFofPzlEU+ngoVB0a7WUHqD3qP53UPP5JAZPMEDNgg6QzGtqH3KKboXZc
D6NliASGzoyTU3ZYgqp0OG5nQFvriyPjYCH+xNXeqVBLVY36VRdV3lPMVeDizG8M
p4qHnylHT6q2tGFGCTh/21P7K91Uvqeyo+Kgpt89kKj+wxCJdSz+wxX5QaRHvGPD
liFAKxuRdVadbielaSCEH1iVnqr0CDLT522yH5zUhUQTvPWWESzS6q+GPRezUD6e
IVPERZWJMIt6/XzDjPPU9jowG0woQI6xTuAxFkX7d6ZkR71nb0truIlnDBRhd4Vs
XO2+seHZ6QnxMuxkFlqxjf1GbzBmiyOPc4vVZe2JXdXtzj2air6Lw9x9gcTfBaPl
pQunGrXFGdLn8HyEiT1cyZ6xNxKTKPOyJ/uiWvMGvvBUCYsnbq6TfjZSqC605m55
Jjyp7vvS9tJKX5/ZddHSAc6NU4aJ1mhaX0XuHeSrYmoFhnLuCBOHk0i6huzAkuRs
zJNBqCW3f9rj4B9Hh88FnJwseHESF+AAErvpm0plvRZJ59hxyQ6LHN2deInzFWLi
weEnECw4B7rUlm2AeaNe3ZuMQIrt0XSOxkqc+ZGxcN+KJbCan3LStPo76r5aIwif
W/kyS7fwMgScWcWHyCOkHllqWHZZu+sUXbgTa8iAxaTZDpMEghZUTOH4JuHEbjkh
/lPfYPINysblYFqmAjJKhokxp8QVrvXUo/NsD67HAtMS5QSNejGJBPDTc+SMytCA
lwZ9iQIrQWFue+95XY0E9hbcA6V5rfoP/z2kVlBTwH9ZQVUFzKqcajaJK9AOoCzo
SPwFQZIiUxdWo9F2ipOCOIE0guDyhpfPOX5UJNMioouvc56yCt8LiK0+nIbyNjWB
OpyeCuHhCSUkhbILRXJdm7m4oa/j+ljwToauclilejGq+CdD7gEveLfvw6htK9bH
urfLisruS9SrDCkQa8sHJ1ECquvswbCaXHpqcTTjxNgRjlvBHfAprB3aspYqzqAq
ozftLiDxzv/Dg63leSrR7GdL4n4dpkm6uoyqaiBX4QIcPAbhL8p0D91GFpFfNv+Y
jr1jzE2H1km4sMvTCkmgRUJNt/m762sH5vCUloTYkUJyzstiaLlTCOW3ge//xtP5
H5qHrwZfSNzd6E1wzFFRHYTmX+yMCcfZPUaH+Z73SQOLCF6VVr8pAo6gX+1W/DaJ
auqbmDO3W2+gVpu3bi+Zs8bG6bBZ2pGolrEOXnThGV/vuHDnOcTqYGSp09Ygjq6k
ZMYWeYeVW4AKW/7nZ6mkN7O+5HZ4R9x5RrpnO632WiFXS0GJFnL+8iSPOoIz4oPe
zUefwKaRgcPrx3J7vqb7IwFPsGsRWUNtnGG3MDA8VaJDNLjYYxuF2487owADCGmQ
VRB06QHvWayKhITHPZt/zoLMrfnelMSbKnTyHPuw7ExB97jL1i8bFHO5HtqkoWE7
z8gyWjoHZ5+T0EvSM8cuGl9q4OGaUD8YzuFfpPWXVdTSgEkeBNl51FJNSrm4xcwb
rvP6NvHz016s+hqwlWk85SIg0EMUKp14Bxz/meQdsj5ORIPOHwc7dJ7s0LORFw5S
/J1Z+IioZHuO4KSjcr4FGzBz3lv/h9eINoXzkap8fhNkIYuFRKrg6UXlainW9gQg
Bx+NGPN+KPye+Nx3aBmBdWDH+ebJThP2toYBxO8Y62m/+IEP+lTSN/RSUTFtxfWz
la8wqCg44e9cppRpk3LEZ13W5PkQdlCdyGakq+a7EsiKujJdGJnfk6afaVPw655d
TBWnHKW/vXFbff9Ac51c/cNzOKtU4pPzgw6jp8wGrS9ouCnuKyVMBId1V+R1Es3B
WLo1OlS//hLLzil3dEtElTiyiah+66Uwh+Pn4M4MqrKqb/C9pIEdkxDfrm4dmfWt
i1PK5fpDwWNOt2nu8juZs7nWUDxDC97H25Rznt527Vw3robIetQqsYEgZdKWBLJc
vu4j7VedxSsnKVQtNc3Vg77m3AjtuBSTnnI0xfT0w8AJnjeQgd7FZ2GPkiJJgZOU
9Rb9r/BhF5zP/1WTybiVrs3/0367qxX7peHO5doVFNvxHJX7tcUtJWxuYmZdh5gh
mRxYDDLG8I0kXMaGRqznQLeCcdkg4iO4ELtxwrRmz3AyKyX56IB8HToPTLEjPJbU
WVKhUhYoKWvnhrCbA9pYqpNbCnFpNesh0ZzdmT5DsHaEp/WLbNKXIlJ8cRcivuPg
sVAbV8PbUSqPgLTR/Kz0LdDdqkHXusaOYF6hTGW3zAqInvmLWwsL3ZwSjbkiPucA
MOnMKu8v0D6n4AQGCq6JHPid33xTaNjzRzo0mAUTzamz9TSLUpbzGKGb+QrtuIA3
JOZjYJTBC/1T571mlSv3H0GO74nZWzZj/tzgLEt46oFdH3MA4iujmts813InxAra
gYPswdNMLdLcKXXaVfdPyvFS5UB2Z+b4+dVx49XFZsaXnRPOgKaAcFpK71Vjye8P
7njleyEs0QBoonhfpQtiOG35l1jDRk36JGHXwLdzM22er2iGJGcn4qDyLf19KHSu
545RVOktJopIVpXW7uUX8X/PUyODw203cNXCA1/7Gk8yvTaBdS9aZKcoMKURG/ZY
jkrcnfbLGt2JaDmHcDnPj940UZGaNULqgdyGXVWNivLfukwIZyS+PyeRIXaqPtCS
YnFP8PSr39zdlHYjh57tDqFW7UE9hVs3IPdwVNY6GQIzAwinBY7U8le4v7+NT6uJ
1YQvRgCBE1DLOL4WUHuyD62UQY/taT4suCgm9fsCtRahxOVZnfJCFYeR/VIwsAXQ
cZaNfzqHr5oR+oDOxfdbn/JwLxzrudrRwhtLtUBhl3vF0v8XZbhyM0kTMw6vYijd
TOQ9D7HI8Yxta0DVKWBPQE03ri76tqOODqxbBXZULGH2HAawJ7qgjSsiyQ1059TD
mFwDOKSopQ+g8TrjZickx5B7TEOTgGsQaGU6FFFCfpgCp5A6ekoERK2H3yTUEo6u
YMdt+HBKxLenrPM2CyITksLl7ZHD4ZeMJIuiAbq0sXNeaJsA/UqV2w3c7d2MmftE
SIdpLm/VxXha+HM2BViBGd0lb+ZW8o+5JNmRBnjAjBopy1YJeLsjbdxfcwiArefw
75By1OlxtO/GnxlTfNMbcg4OwBn6h2QMsJQGssr32hNFX02wsKRUWRL++h7oxapY
TzRJx13EZqxtljE+ZQLXypjSr2x3F+6dlz8FVemd5ypDQXVrLJqLPG04bB1BI62i
ASgY5F+JQu2RTDklzPDIas2ueVTGtpSXQnrREWVX1ieDn/GxVI2pOm82up141AP8
QikymWg1KolrPMeECa6ZqNLFKVGvfjqf6iCphlatEMQ6Z80xuqQcN2Su2wyFqvv8
qgf6RR73wWidX59Ja+k9hD6EXkiu4NB1ic9dTKidYaRxkvxJaA9DMxd3gNafTZld
p11qbuetJ+LlyjMhacOzXYZtMCP2XzBf6JIXnmen10vcL/vKgNPot8KISN+ChkN1
CbeoDJTqJJVZAdfPtkFplW1TFZgNDv2SB7efJod4uRkLbF7fhPIGgo5QVInhDsvB
sE0GpHJnIET5F39c0tubu3XcbQYU675vxiS8zA64gAIaNU961ONLJf10kbbFjdYV
Q9R5U05C6iLhw1ey+UJoVTBxYtFnov0N2SLBvkzryAsl/xemG5JDS9FiSXML9mUJ
ajFH8oTvXFD7dSWPPThTAF5UssjELhCpdOTPprpu9wS1+8q+RBzs3N8XbSgiCjBL
pLhFgjnHecPQuk73lDHmcRIYlrk13K3aIlwkIodQqyASqAAXuq6idT7ajfsLIgwg
ncVJQ1YSyKvQEcxzhdUnBz0Rxb+bRBujP76Kw2JvCqB4fAcS/ConhK0Ewft7Bg2g
EBCTXFGXlcQSisoAgbMvYwuWiBAeDTJGVw0O8yoQ+v34Sj6B2Pt3kJsc/h5vpoQU
F+qemZ9XgqcWYOzIm9hZ/aAKtIb0fBy1WhWg8njRTwXIN9ak4nMLFNUJ5AHKHciD
MOrrE6eusSHcsG7xf925ViVBacx6iKj8UtdEp0VNA6zpRobZBDUCTiP44cHR6qiT
V8wFMJ0Owc/fn/j9EV2ayXtwF2xYxOlX7OG/IftCTZy0kAaubGUSD6s3F8qkvtg0
SpWw60wJkg+ENfajZ0zeIOIWFORfG0SEioj6WQKxbUbVdhxeOewwk5RF2xdyqBzh
T2REtf0rQSObB7D8sBzFVwkVdi5STHeexZbBfPpWYe4JBqoSF9NIhNF6CFtty1K9
ZcXRCa3MmsxacO/YRwxnhohr/MksB0mNvnJTC9u+D0dqahjDC8gDlayxPK1BWCxI
fdb8wT24Xd4UW3c78i1iF3z2xW/FxZCPJ7ttyNVZwkLb7PuctzOBuJMWDPZzLX1c
TF4Nt5WgNYzrCQqR/uiH38YzlNueySqHD416J1V4he61ODEzv8jFAA2yrkzMf2nw
svi8sfj42FbzykBcMvI1zNXsnodCJGP3GUVGPoLR8o8RdvIqQ9nlTBcNc5LXuyMH
u8WtJ0STYmihjr8oY7MV9MK4mGt/bL4xjIs93rc3cqL7sltfZy2lG9UGFFuar95T
Qh9vpxz65Tr/Zu97ovLWZtyx7iHrbJdeottNiiaZ7NzPJNL1uGPpaxYylwCH7y55
3Oe8ic4sS7EigvYzaJLA7ZrUDlMNgsDVlc8KUp1sCZuP4pEpXSdhkNOcREFRZ8W8
LZETi5ogTcGxKd1XolqzwS4mGPBcLabU3d+rHrwv3mNO781VfNh/tFnQV4guSwNX
4rYkEqR4deIt6PepN5oYX3xZ+07yfrKSkyvSf5E02oT8xlX7M93pIIHZQ3klXs+N
NLGjPKLj24zD95cCjujf/S2ei/TJoUYH5L7t5FHPMPwNzNUx2y404PmZtjMLPtIb
kPkNOhbgjbd/37P8oUH3hVQjYsG+phDa85L4IaB54EE2/LUZybD05AP4LFIb6mDc
gMgXeeoR+pLQsqZiKQIctTeF75BZ/dm4R0+NIEtvxpWNNHolFNV5dWFgA7jkE7i0
Bg6HFVj8aT/M1b+P4GhEHEMEnBeB1h1ixf7Tu++5Wv9+UR6rLsTQBwU32T0NZSKw
8qB9pqmUDvZHQlqxPZGv8EDslF7bfRh8h1jgZmZGZlupxdU2yXq7N4Q7MK+aQlFC
a/8A0RMZ7dXb/AJgDsGgAMH3QHaZ99S543HoNyWt5hFDpMn40o7NbnljuOavXong
B5Hyz1fhPMUfgsS02hwRSqdvNQDm4uS3NRhDfvPBXEDmAALOAg5b8LfbzhOdwO2p
SRFPH2U0UwDlzOZBPChfLWMJC7EQNwWGYh+/rDJMFujXMSYlVACs1jSomaKOU+or
B2ZCstOkx4EozVmcR57A0C6hcbMZzpfqSFVOv+Oz6cxm0PX+9xi3w8XQ/Qev8NMt
dQrjC753asou5jk9uv8vGpCLQVhcVpnOexZiwOlHKmIQXR6K5USyPQzCWF1l1v1m
uvYibKztip/jMyNApdcU49o6AnIBPIC/0gh+KsNIxeJXLpgLNA5sj3iujsGCZ/Fg
AjkqnSAPq613FzVw+MJDOqDGdOCloNu/FEykWutEjwGl9u7/I0zJOIT4in4/cVu/
RFFNVrDQBFcvG1f6jpX85gPo9aFIaouQWTd0fuhf1WLjdRUMnMV2NzrBYz0nn+UV
iYtCcqPqyR3/QW7ynhM+rLXR0qzwZHz4J+fkVIqbfifz0bW+oqhRfJk4BBqFp+1V
PZSlpvrjuu5iJ9CEtVWA/YVX0fxFOpmb/sFJ1xdx7apYtX0GSSfeyLzivAiVJhsP
Q/muCCk3IfjrK5tL70JeoDUlPosvIFRoNqU9UKwxN22igS7xv6sucYdA4cebAxGd
Qlcj6cb8f9pV9/vdSnOTbr6WrCxUAcKF+T3vhuWna/2+N9ItOQsK4K3cD8R0+scE
XiCeL5IITkiYm/7Ss41hNCxOmyZN9G2QeKMkz3OhFcT7//fcfnvEjZG7Cs3uIzr8
9Co70/jr9D0uCADF0MKVUKYxeMdY28pn1EBe+TneBmgFsIaLuHlQ8qjI+QPtVVqa
TEtfp+CW+0q5pMRrDcKcORx5oVTB9//DnP/ecwFtwnJ0Pxz6/ED3XAIKGRn5XwSo
7qrECATIgUEDWzAEdeG63o1ab2bbq2MvIaB/cf2Bw9QZqJrtV627Q32w2f93khOf
fBz054szuQ4riZOMrqkn02RXuNU7U4/ZUFyIPBtCmei05n6lF78txGwMdNYNu5sn
WZrnHQY98Mptd8Vg8MRmvZT5cQQrWAFAEGN6OyEizrpFZKYyi/oz96bvLh0ZXIW1
Aj0gbcar+Gsj5DzMZhv3jeYcDVGl4a7SjOMGudSweOd00LU0A0e6pnQBJhFUwqVK
n7ekcnnfz1EKyK83lM+ZrEQOUNPo1KbV0nVaq1du7+9SKAtkQL9jnmucQ5iSyMnu
/Sfujjf8B1DkXcokJCbMvDKUtb/EJ3Ch/Trph5nQ4G98toq2afDB7DPsVRTs0or4
acI9O2IYcTf8J8hQJl7Rx7+ov2zIfCU4O/vhJH/MXjWLuA1JcaNK2i9gR05QrMtT
pCCTEVUoOP74aHjmeqYZRfeapr6EIUz+r0cKgv0ql2y1CIuJ8taop28uv+7R3HJv
4a069ev5DkSMD1Oy3uOFmkXwrLUD1Q1dPAZWbWMXJGEGGKq+aao2loaS1amG5VUF
l8wdn+YfCW7V+C3/g3gaNlq+RyDzOxPUoxqeYknqzsDm60z99+alRcTUefV/EqTr
ymX2hFGiyZPZyV/n8bMtVQXiHIq4Hl3oqHBztxezyJ6ouBUJwz9Uy7wEvOX6aGM+
C9yRX5cDndtv6pA3dONmjhCcVVoQADLqwiN3hEB1KWhJ2flBcL1b/rLEh9deJ5qx
EBg5rrE+SPTbzlsUeQhkJY/paQQ2ponRcoKXBcn1TS0lcS6LQkmWKpFhRwUuiBJP
28kucENIqAT4ns5W70LFjJwoTv7KeWjk+YvfRWqVBMuHmQDTuHyH871HjYzDidv4
hK2p7JNk/lGz+s+kJE/gcKuvpHttnx/Skv7DY3qgPpg+5JBeV9TGSih8d1ZSS3YF
gUj2XVr/QmLFNuTQA1pDvE5FujdtvRsSN0Ek9ELZepiAc1uPkgGhIYkTnBzfy5Zk
y5dzmG50ZpKMzswymSxJqC1y6lEU2W4o3Pnhw31FJuPPE82c8SWwdNG/9MTh3mcR
pWGQzMqJEAwjp77mZNmkIvHXMyLVQ+2yUk4ILDnJ45e9fs3UDbDJlJ+JxtuLYgx0
txVzHaWSO04+LzlcEB+c9n67pLTcE4XtGStbkKyb25wzjrEaM/jNoRu90tVLpeGZ
Np33VEdMskGUVs2ntwXTrKgmjAxL1+umnCTYAcpxB4LppOW+PCvRChnFgRL+BwNj
A76JJX2QWXR66qR1FeZhT6upvcIsn9tbxyffQlGv/iqhYuejrP6qkM/hvaxXx7ma
c1wQ4nRdULaWQ54Jq+T9OS9bK2WzqXHwksOnl1Cku6BkUT2jW3CppdCiNP5Z1p4v
0b74zrdcNY9FQJQ0ihdfDHediGUBdTCqyVwe6SS/66mNe0NN5SpU3Nt3nf6vmp5f
TMuTfzfkClYjJ9HQsuQSyVSpuKLEp/lKydr7CUqnVc+MWkfj8F2DTd56FiH5WCrd
C+RYaiPHjBFwdKHQU6wKW9zV7HTzRPI6UOGMf1Jpi7oiucfrrTvGqB/9X6dUatwx
0vA3UV2C3THxtlm8KL9z1l7jiGh6u65Y+3cEdkIHx3jMz1qgZTDZ6JmqzYlqHhvP
kLAAB9PnLzcljOAQ3HYDAql5O2d4WYAdOhmuDJkfKRgEN2H2wBA5zMh4mj4ihHBo
6BRgR5u2Ayzr7RPvywPZdmSFCt2gkh27oKlBvLuHfnQkYhfsaO6LAt4TZaK6TJsH
mucomRVorBuyTCnYNrUKL2/a9iawz5DlVF0nGKxYUM5GmwxlFVk5pBTbdqhNolj3
EA+juJ8kjADAS9LBDQ6E4/3Tm9agS1pj+UH3hzU54c7JWrmMaRK9aoJ45hmeik6t
FR/Jxp7SdAngOFvf6B461F6K6hZPVaq7dCDqn0n7tuuMRcOIR1mV0xM4dlW7qHmy
H4kCZIjAG4KvXAdK9glTuV+iAEWt57u5P4UBwCVB33vo2CFquABpypK/YDDmsdfl
Vuzy2Xu0bbAbxYA7f1eJA98qbynY6Iipr93/t9/enifzyVHsS/xSWGDNcr+wlNjT
O6PoaN/8UZql0PZZpxmRjw1XP5JfVqmg7zlVcVLqZwPdmLO1tMafJoGbAjuZq0gj
Qa5b2ZyhHrYlqYeZEp6UzBo4mQOxTs/UCj+o8AcpVjdOPr4vS+L7t7ZJHUoRAN4s
5DzPRlt4u/6NePoVfNgwHZVLf14siX4kvST2Afk6zm5YSQ+7nsXguY+qzH9f1Mf/
C78qfi+muQJu1gFhkrQCq1/27siN3+NCdt7pgPJzwXc+kAX7k6j3Qdfntn0HY7zC
kTdQWJ4n7giRXRYKrlJAPjxoLDxZ1YJMMWqmDl1LNvyQa3wy4OjNO1IBCQqRmljM
vrIjU4F/+PXrK1fMO4B6MrYEHCkLlzlHm01mT31muuebCW7s8nbBUU1fjbS9ndt7
kwip9gh8lba6BdVHKFrTzwivnkcfrmrMhyfztHmzAuRXYPo1sf0YQsERlmEoWF3O
aGrhmD+dcwbnLYRZ83JA8jCey8VB9u/8C8AW1r5pA6SL9zaCRXQEB6r+BvY9xwEi
dScWMnwKE0LzE1QJEfUhYjPrUPXB/FVH8hdsh1qPbXkNXjPwcMgGDr0xaw8RydJa
xmfpClOh8CmMBooRMFoQ6qVS34pN60XApYtzAQiSzL8QhMg8lBlkHpTrL97HE9dM
D/QTKQH8d7ePg706coJvQ102mMmcOnJHyrbUkMgjTpG3vosHgsTArsfJw0wpQWb1
Q4Vf/M6uMTpWA9hg8smQjraxwua0VCQzD+WzpgnS5KS66bmbNhT6NDHaqaUJ57K3
WJRwgFm9qUtHvKHRwGajLNubKZo1ubruEo79ZCZkLXwgpDE7vQPKNh6vTbNQqiRl
UTXOJ0f5CWjKVQzU3Gy5Du2vZmglISeS6nCvhjsDB+BI30NkCAmd1mbiA0HepKqo
nYVlydJtAtTsk/dgI37PgerGBQrAU1e4BctCPk59hFHrxwlqdmoCvAKt/r3S1KWu
MPko59YNIQjR2pPZ5Q/T4R7j3h+OhZUPsb6Qk1cIDhmO9R/FS8LxmIGdhXY3I6jl
/sjxehrkx1ePIj3KmWG683tJZhuTKKjkQFPKZSeb/JIQTnvbWp/0sat0yEYeBT5/
6phzNUjARAgMYQkE+iMNtjBppd0R2Wm5ElFVL07KROWJy6ZHnRP9+AaqfY5n8s71
GTpc/ZyPBvANXLKuOZWzN32jlh38KKCje+LY6gqZclw9tvdBG6nH7kYz2plOJg5q
1E5w8T7cK6/2Us8iTM13M+cs56J+zCW60NM8rIrQr/Xg4Sfze++AIIO98B2IIqvG
/OvuuJKvLyidlPe4RalIh63FnC4AxVTzhNaIVU2Q3SK7kUcXMM4rQsFBHwbBZKBU
n2Rx9uuwVHX8wHIvXLt+KHacQTIli2cbobNmmCp234uG/IkjlF0KMCC9B41tSGuI
xxqmoLDQOBEBCbs1sDegQT0XumCQ4qrIFG2YvWq3UvjxuLX+LSxaRWvKfQ1/FKUc
+8MBTqRH7ewDJ5seULJV5U8cf/0bMEzB9q6MUTovGRaE8516QEty01Gjpt/hD3ns
TCeg746XaoA2C0CEP8RKv3+KLy2srMkjGB+kFPkkovZUHBLhn8/VTOl5YsvlO1VU
j38MZtUFtZyHbcu3QcZcVxCI7lJEL7LS1sNqyIWS9DIM3E9VrMEyklXG9xcrVGG/
ertnSIVr4Yn6X4r4dXnALlsABCI1kLszf3HGYxz5xdSobvVwU0BU4cO/KP6qs9NF
JnWuPLvQEhlmtHot61w6OpaO3Ho/V+9BnfNJisj3KrNFV/V/GjGLc8az26aH4S+2
tDdhs1fQKj/3dygbV8YJ6M1eEy4cs0rQ3N5vSM/U6VAZw5aCnj0djky7CgL+M9lK
efbkZpzdyrJTSq/Y3twETr3xDLTS/6rRGRC2buL3YVxxPjbtxW0U5PF3ob3GOC9J
OvzPoMxMg/KHORuegjbqbLxvZ1kJlmCq2pNWplPznHzz12kE+y0MAsZbpcpgshgQ
+FvkLRHBKHEegZx+VHJwrQI8/aQMQ1H3Rj2hUZV78/VchtnOwTcABVINZWYuzsjD
V9CYS70jkOmwyjEJ60HOZuRV0KKP7+jNZwnLxgmq1Kk8WLPDvS5H6vrE77AKTUdp
31JHGCb40nXERfLdzj7KIIBp+ajpbp+5/spnaicdUT0M3WQ7We6xfIFtMwcbN6Jp
Z633ba/X+l0Yj/oi3PGL89HwNDKm97o3+2cLazQECTSypLNp+dH/8ZtQ4P0QEAMP
9+xsht5lvCyWxkYOFZaSdulP6xw6zaMB38StkQ0yWz1Vpb3zg/82fXVzEfl60U0a
gZecg514OoVA+X9DNGaEq9tXy+Ldb/YyjB0EJXicnKrTX/I+HnZBalwsEvr3uveo
aD91yqzQGCV4KOXj0KhH9INBG8FV2m5O/EqOqgrlq5pC7zyDpOLmxve3SKEuVRBZ
mwRefn/F04ELuBbHfynRDBSpqO9dy9k+ytJ+rhwRug+X2mt+mJiP0dI+w8akjRzk
gSW5ycrqq/vfG6rhD+Lv6Byz2I01nKAy+XUJWeXIES36+vJajHHRGp3bh9ufolud
cZ5VRjNAOXRqNsxhN9Ag4lbGfrEOIBN0Oz8eS479b0J2YQzgPdWbJREIW/QcxxXZ
UoGkvqXUlP0jFnpjtMh8UP82gbMFnlBbyqgxMFF1VVMIhAq7fy1l0xZ8VqCs+Zsw
wwUiGUNyRZINWW+exohzx3+xxIiXvm9wKU9L3mm3ERtDDhsPsDGQND5d8gq+aEkt
x+0JflDY4ZLC/OsxN+LR/colcwQZJjEjCVLJlBtKnoYbyPixOpjvXykgN8pC7w49
xf2hgpHNWMfDooxzDV75exTsCZGM/4wkvH0Cq18h2EgsbIOB/q2FWRqXItreQn0M
KPxAJLPifjIeRfX3556iz0jopkWuL7NLw80VcJiiTIKUCiR7YFOig91OiNmdi9sP
01dliAJSuiwIDb0dYRmH/eyFtjldVNZ1MM5m6REODTGFJCedShVKIJra6iX1dBkE
E+GsWwo3r+iN55lL7mLcyoGN4bC6FwZDsItd9IjimmsDB1Ug03exhnnmogEGVz5M
y1wmNXpQ7qlfgwRQn+iS99cO9rgtQtmZCJrqph6BNybRKTmyi/HxXxHo8nXQ0I65
3NhbzGLX555RWXkEltqisM6TiAMuWxLnGIzf6+n71qmOdrKGxdZ1rmu3iFSjDvMg
rD3H4TJQx7T3mw6CChB63PKo3AekNVdXqWAG4cGhcf7lhrcFKZ7soSiM3xYyVHKW
TL7svkM8j1LGaL3IclV/j9Pv1Va3bLJC+KM6piaRuSBBqXkAx8ZyIwWm9lP2b4rV
ukRrZeCJAYb5x0nsC9UWjQ9y0+L9W8Qr1SytQBftTMWXTrZFUJemvYqWDadzTqAU
qQqdtkRELnJ8D7/E9pGFGsfxSzYlcoGnULGunGGd1oSzgK8FLlfo8y489hAwIrKT
tp0VS6HF2mC/8WJu2+j9BQ5PHbuFa3Rdhpbj5CpxcdY/EpwmW726C5xK2EE8tzHP
PJSI9oU1SPzLuIvkzFXP7t/0rFG3WVXcMIFVXxoPGXgs8udEhU8UOIGNcYH23pXH
XJvLxr0u6uPRrj9jW800AQ2rxelXsBeHLihegSNb3+H25QsRtFF7cdNedjDaRE7B
/PRz+jroIPbkD3I+QgTr3zQFsaUDmvmRE5bZyJbTB5Qk+NAQfltskgk7ppUUvuQq
Iv3V5UAJC0XQQFRcqLyuPGWh0ahNmJmJ9nVN5JST18YE9H/taMiIso3ocnihTITj
DuSF5cXrQmWDe9n5G3hlm5Sgm5rIFTC3j8yP/QPEQao+wvbpKXVZKa1YaaYZkDIA
CAFvgXw/nVCh5OjPnmLFRITgaOtslTMXehOJPxa7w1NiMnw/+uOw6O1zjFWLu8KP
t8bc4n4RpRO3+XqP+GjD6fuY8Q5Hq5kxe3WTzBQLj746sap4ky5y4gavx/k1IxP2
pVmfTtPXwCP3l97GXKxd4wDtroCfekJnXAy77vs706BCSS2ij30Y6mV9WePZWDa/
oHdCq2GGbt7I/0L1Ys+zaTSxZHuSIx24cRfEmF5XDbdi9TmnGQFHXIXAAshv3ZsB
qU7LmDEYxOquDvZrCWXvzTJ2LAoD5QanAFgwZCJ8riiyq2uVNOnKTwPKsSPv0Q1t
biruwyVgu+B1p5JwbHykbLC9jNpE8SKHCfyZs1Bz7dwJoTrPWGeYyDu9N0utIg+6
wgpH2uPnsosDCZ4nfk9ktYHdcYgTG8foGxyXz28g9CDev4FiIq5SgDGKh7JrI/jY
9/S58O72hMlA1smH7ZHg01iKF2XrGtMcPAZkZcxRYl9MBM8BtH0QVHx/Ec73VGOH
MOJLphAd7+l2z36NY5KNMuZ1DQzjlwi5nqp19qz8xtmu3aHoy4W6skFZQHaj5Pc8
6mZF5zQiqiDDHG3bQoUtyawYK8iVAZoRfoBdrsI2GBrf6Uhj5XUbumSd4YlRMjN5
7nUbqnZBlhrbiyl8w28XtjQsVHwIk/4rmqQg/Joru43nZo8jV8iBL3rsvQwrzhQd
6nI8+oIQSKsjOyv5gGWHL9ZpZu+tG3w62Icv+A+kxMjExCY0NCLdyOcjPcwNRaad
VFvx70lJ99f8VYggVGY4GY25y7sw07VKF0ebUOKgWwVVjZ4YwZy2a4d0PrSeJlTm
QgBlS3C99riE+Jgu+7gjiBLxNDbutmVoH4Ar6KMZi/6ZLTEUehe6zilVwuNMc7rv
U6sSD6ox/Cuj0Y9kJ40KJpaEmRZkImPO04WTAzigq9iIBG032DbJOFOr/DR7CWyf
fWiEaxa3p179O+b4FAvVGSO7j2s9oxx01jbrpbM9/0JzL3AKM5OWJF7ZNcLlBadV
JuAY4OmiUVntfaQV14kEPWqBpjatkRu37SpnrT/QwuhBP0ld1Acz2y+kJhjpXyxb
4CuInljPSwbkU8IJ/94ddAb/BBYDy5kWgKzlN80bZ9ZKf3UMwK0kJ+tnny7uNRb5
iyvXSq2fGYUfkc39X0otCbm1V0Ibu0gF9b+bu/zhRYERdKQiYcPFhmDAPxICcLQK
KBmx12bQDye5sc3q0pDuTGvMmP9njmbzRec6i/i0yJrS+n6Sav5mypK6GGYU9hfL
u3Y/vQJSMQ5Zl/FGwd6aVGM22//8n+KcvUS7eCKjN2PFr4XfdfELC31NXDl7wvSu
utep0lSizjMgcqQVr6y6QxQxDvhRPahudrIASRq60r/rhGcVPFRu9A+PzYIuNuXP
Wj4reAup8kJb6Tr7TVPO+ZBUjGpMBhJRcRsqBGGOAOR8vML+OTt0bb9bzZ8OVHI7
jNe9LC68BNQY0MoMYai+wPFgrWh+g4RvpmgthLhRC8n/DVWIE32t/wFHQEC3kG6W
u2bvc8i88Prd0y6iG9QTgLx5m4xFc3FrWqfhJaSYPR6oa+6f2nOCkJmg+ggIyQFf
xz9SALUOliNphAVWta/Z6q+e3rPJD/UhxaVegDdVUrPojmmf33wQotH77Lk0Rx4X
QHUY+ClmNXlHtPVO6sIPHb54wZEy4pKaK+a9BRQb0J3nI4Mfk2R3yvrIZVqqYD7t
yFMvv2BLxKxHpmgsWLadS/G22mQxHbkQCdKfTnCfizQy3BLwy7OiV/ZTcuaE3nC2
DzHUmfitj0oPdA1qn6PTQivDqupqQZolcquGIEBQHt6rmOCgJ7hYvETuaIb6EnTN
S6V/1c5fcyNuq1GjpItZ9szV9J8zbwwgFS0fRv5vHBCkhs969B9A8ftjHvJZ1h0Z
0zNXjT1N3F3NYo5FfXIueTW5L1G1OIE9Hx+tEnO70Gq2DDEhepAr9aQS6sp3ITvL
GFLY8bCBTPGMNIBz5HcioGf8Ut/rlQf8Ub0WY+7Ge8ka2fGPUI5enZFH9rFGldjU
gyNkCBAshjL0aKkF2LzvhmIHQIgOgeNIwD6zZP1Fm1nK7azSQudpzb7xogfPUBDj
rfD9sBUstRyaiM28veRlMSPDj4ffg8e5/AuQoPq6V09AvImUXdadzXNlgSl1Roww
E9K1X7Ir7yyBjJfNmZLGP5X4Ytb6MO+Ze57xcBuG796R/Jspu4bIt4A7H8kWnbJq
sBiYhPDzOPTLbffjWx0t8ge6Md7xSeIkLYSfshnySKJUhpt+guRlQAPGdz8MSqUZ
UkXcm4PULQHaQfq7GBTwE9aTpp/bC5RdeS57sbYjDDpHONY8MZE9w/6WepxSZPgu
Hr+ekw5+0WfxS/0gXfNjjX0PobxG2M7vcmtRPLODvrJbsIWoS+SGKXq4VepSSI33
pSc716ZLQchEj1c9kBtlOa5019LzHieJ5H9rXTM7ngbQFAuiZrrEOA4AyZF6Srlc
VEi5gTDJKRZZUjXRg9yW0Kffdw/qQJBmQ/2y7JEGpmhLZ2/eQJ0+Il8f+8eWwS+8
iSsL+Fdk+lBFQMnzE3T/4pOr2/NwkssSnbM7vKwGQbcWzhjydYwYh93eZcaMCG8v
UIMbnRIrv7SVrdQ3pU2JdXahDSGVLTz33P8m+VDaHmr3cIYSBHWWOrXfhB0OG6Yp
M37dYKn/j5c5IUO2OOAIeYQ0iWeJSAkMnr77ANdQ5GxGR1c1ZBURhky/p/dJmkNT
hQP1bufW9u40Nz9EkDGCV1nHQjun46hAcoS5g4IA1iB1Hut0ENb7Ayb+wxlOKeAZ
bLcKSvHy3hsN5KF8XCTho4veIBrMUZCf+0d+FJ3HO2fc4n5CWgbqAeYHWDcWeBkU
Oe5DiesQ97TEr9j+xdTe5FA3XOPBlOEGy5X8lr55RNZNS33gOul8/1FHuGqMi/92
p6YIQFhyH3ACHBbSNEAnOxJqbkiQS3mHVBeSVJH/LWN6fyRz4+74WoUp1ywnSdDh
6hBDDotZDxFLLLoZFLJ1zPcVFBv9+FbS5qBR1Y991pH9rKKZaiWZ0YXJFpLfa2Nd
Wv1UqSeN6kHNn+C9EFJflnKX3BgZOrLmsEnwGCbPxLVHbak/9Q3Z1oGsh46uvqHT
fJ7j4HIjT5ImjnCQoe0BUXgVg3VGUMJr/SyiU2CZtv5NwJPIS0Z9wGLUncffAwkX
RxDYAUtBSTWzx32/ejlQnAhVf9stHghQCIuxBr1nFJ3beiDsvThawxMKQEyvqNCh
blgAvLyD/BwGowJrZ0AdZNJp8J3b+kDQYwl5dxAfnYI+GewIGxY1M3m5+KpSH9C9
ekERk4Tc3bWSh7tI9t+y9M56KN4DE4mRJxYvKJ8AhOzUuwWsCdwEh6OLcJSWlHaQ
c5rfQUh14yX3jRbBDNto2fi/23S4SAJl4HFOu9gisrRcdyJbNDoAz8eGuk4PkkN6
nMtwp5F4y8Infg3fGKdHXKcR63IZtMg6mg6LuP9ck4v82ZXWbta/8IEKIDo+X9tt
AtbTbO//20Sb8mQa/ptsAscNEUWNqZiOHZE9itag1dPvoG0k4oafSf7QuH2R7Bo7
qB6vWibQQZe+ZHIwdXZuX56K0WjbCS+miooZjt0ZlqBLysE3ipkNUX8OQ1vc98Zo
Al8hvioe0f273KsMxuw4RzUZ4puv6vphv1abz+6HT14QZVWWnp3TJWkdEwxiBUog
tk2M/i9ecZTjh7z6Zwo0PEj3PYRx6h3V3XDBq398BeBsVV/mrReLBFT7v2GYvk/d
BroCz7Dc+YdQRMs/79L+8AP6f7/gKRQoFdpx0qN5S/Mw+bk4yg5sxg6pkZ139j9I
Fp5GJqaw1zUVqAGl8Hifxxwko7vcIvn/AqV9da4Ytt3h9QnZKOTtKjroq0GE36C2
9cCTGeDzIu3zEhgt4gvr4+GI0AFs6dt7gNP8YpziEQav/nknZQyn3W+l99rhXI8u
Kfk6w5dkhy0VhijCZY7pu/riA/Q31T92He3qhkUUrVz7xBQt9fJ83/2Mz0wHqEID
lPnWi1gIJuNJ1XL8ict9Lc43lRUgZfQwbiXs6Sn/c35O0RBISOAyeszVKheIUjZ2
HkAglzcHWk5ecn+X621d27JrUN4+IEI6Q0uoYFKqav070ka920/LbG7Arrfq12R+
57t+U8MiZD2pTqonI6803H3SxWqSuMsRF3T2RQxAcAzs3p8VqplhZWvUKFz5G7fq
TOjsa/g73dEJgWKOw/gEJEGrbkH6tO5Wb67vsFjGH9PAnkXYfb6Fgix4DnCzk1Qs
npLTihYb+yEKPpF04lrtK092+Kkckcy5u1FlqMZjJvRVbOYU6IO6w8MI6zB8Mdz3
W7MC0KeKN6DSPQHhUAPLDvAHt2DEVF/b0eh9gaPtEacEf3IDtVtda4zIsjYK0wz/
pAUXaMDZbhGLa70BtexzY/5/GsWPQBApElHOEyTXl8WSJCQ6FbywjDXFDE+0BMNP
SNskuI4Itc+KrmS6bjd/9gNYoMkOkipPUSqRxYUBhYrkFuirayNajq8Ipxr2Rswe
S8ndizXfc5xYZPu7rPe5eMzHkcqa3PHOuR6I4GPrpdrNisyvX4XJTZfMa0VO5NX2
DpnlHHK5LQmqB+fB8OxuSXs0M5nGpDB1DqnmaRrLkSbRJQiAds2mEnsus/Cu8+rE
BeMPmUe4JBhp51Q4ZgUKlS4yz9oDO2XQaIWeChJotCDIKryK2VlZ5OTuT/j9QOTS
w7g2eUIu0Aopu2/+spk7bGjmMUFSQFKCn5jDU2i6gwmQgmZhj0Se/qsW5NOsb7rw
6dgSfZIWmUCXiH6+QyX6gRAWOMKkPJIJV4fTtgZiwsmYhHFxv97tU4SNbrtmYwVc
fZlzH/bHPF7RvKgmirJF2rxozYCazDQkvTgDPCwKrnzcBun1Z+JGzayeWwAQSmMZ
aQ+ZbAiUuEQxZ8Wuu45RCk62v0/NHLf5fAvHyGAwXE7EmbcAJ/Mbp4lzWkaS4s/8
MPnOPBrdjYeL5N9fuxNaRxVKzM2IxBiek8U1tFTk8eihAzlSUSB0E9dWLVblRnNv
yQubf2+4gm/DN/TeErbigL9oql27gGP8oo5hTFYwVKvf+yt6G4DAHJ/cVVJ697mY
DCg5iW0Tm/0Vy9evU4H0gMRDSfWaURl5d8N71LMqbzd0XxipnhhX/zomL7T71mf+
A+5CgkatDbB50wpGDQ7ZBLL8Hql6KcP8pO4RrYkgEozTIFzc2FRy7o4YRcv1kLp6
HsA2FFRTDA7ECOCECYzF9ey15RXe+hFkOUrX9lyzLzLTaUvz4VFcxSmXdsRusjKx
KqXkSUPZNV3j+ThSuoxR3QmAHI1TYLXqAx0izNvVli8Jms9uSL3PkfQpGa2tQZ2J
k5sd8l91WIZicoE9OYcMCAZsBZzqhhSqHKLhxNj6mJ/fRKySuXcJhOV36yQcXg/C
O6Y2OSukWUafgSKoOP1tQeCmDzD4hEPIerf0Tkjs+S4Lg5KrhDxLA5ALF5+8yA4H
WDVASGUocExw0Y1z1Xx7IQGzYFeD5fE5fXviIsmJQZI0IONLJqNjx9y07ZSlLK71
ZZjeJTX9dv7LcqvH9+QfzOylQVI6o87L5p1Js/gEZURjUD+1LUDWcFsYsCKcxSke
E3q+rEb2mnf9EM1Mvw1beETAsYbkGhGwpBolTj3zqxzOwmL2zKXfubefYvxcjRZA
H4b2pEWddBfOmKe75zC3QL0AazUKvk71q35COiprcvRkSIH92qqHSeiVGT+dfbd6
KRpKqg1+Un/4v+0s7l+GrgjDXhMxMfxFyFvYS41YT0Pz8s6thSY3jaf3THP3XBU4
I/P8FX4vRawxJ/vi7QCMPqqBtqc8pZK2t3/kPxj/Jwk3ZaomVSTE7MPCZbFoVGKQ
FvXB46IK/QiqvbcNOekaptsTvTXnX9PQpiJb0EaYcr8S3jAdO6uZz4uOubcP6PGa
83ELWxmYzw0yl9Hr78bic6c0hOQu2CmBmEsElOvdmjYZ9hXwzKL8d5exdoTmt0Nt
+GHuQN4zvfKaCp3xwi1w7AODpk9bmVUfaflcmTHdD4mBeCGHXQf7vo//0REaZlNE
+ed2088DIhtjV5DGKC8KLF8KYzkhAo96XBRFzVZH0gpwrJzFm201bCM+/hH3nItK
WRn8eCunIjUSbPzgm1jghBqhMwYjFuNnRcFIrIpZ5hL2UUod2CgYDH9xINgiYiR7
+UteXYry+jNY6gKTWiemVx1jUpjvomH1etpO5d7c88BfCJpkPANyhdbVtDhPZoPZ
m6qeRL3bhWkNYdyPywPwcFWB8J5wD2a8C+J8egpg6OlAYzTXIX9LGT3A3clR5/tF
sfPf7CtQfWJ1YZNR/yxb/9dwu1OTT96e9dpKq+TyjbfMd7Ca67QduXyksQZRElK/
qkwx8gkwRt6p7xGdcmVyDgleixU1Pbq+p/H4inADovvHmtgDfh/L6KnahSSPd4PU
q/FS7jav8eWmpyIe+pBhu2ivQL903qFpFMnAmw7H6L4GZB0Mc/wFnhPChaRvdcvK
OBlXcUlUyKc4cBdrlwRDCTAeU4ckeI9BGM7jhe7szMhQ6WN9oQSU7p9cMHTPT56c
akkbwheu7MfwMWtAVIAF4kjLLCQ7K5bGacYm+TV9tFJ8+tKNqGXqJhqRdkyvwxOB
r8/77/J5/upPTVbdnbFcnbxHTrTFZ2tsw44JeG78RWzqnsr+jjWwsTGU7ulS4UJP
+2mxVq68IS6fH/IhMzjXGYJdcs5aE1QXKygwCcXUgycGuXI6BnXnIg599yC4v3qa
n9nRVWaVAGpHQsCgMVQJglEnL6ZRMIvlUKyyOjNsWpp+niPso41Gi6gRZTXXM7Vz
6E7K6JUwtAN0LvyBmifpf0ngEk34V5pREmTLVINKBUnUNxAcokANm5tBkoqsHxlB
/XeTYpk7RbkWixWwk8v7WMO/1xtnRQJ0AyjfwRebiY2hC0bG2kuL9QvPVcoT2KFE
55MWqs6TGH1ap+VL5QafrifUCgwnsvzHZ4KAO/bmQ5RriGaY3lywyj8yaTZZpsud
6EOCTdfDEjhp+a9X8DXkHkrVg8+qCq5DWoIf6S5kMl3oqahL/fH7upTzsiHoY/vM
7Xkr2+U3kAMaQkxZBXbvShzclEQN5wj7lbXcoeD4GVzXQaiyaVWK3eUDmSHTp/pS
7bUbcLAI4UrFdd7ARpw1LqWZVVU18ADtfAJyLjHOFJnr9FXuAD1nAo4mgS3VVBah
HLdD3iZdYkx6WgmzQshyUhelu7tTvIj9fN1XL562zHVzkmhvA8zofRPSiDbuRNxv
o2neNEw0OtCvEmHSdiKlMzXlMRgrg5iJdhkb9C9wySnk4CkCuwg9hwjeVTH0G9h5
qliQxvadvMS8IGzbLhVvEf6qP2m3MR0QACxfI0HiLaPBDDQlryY0b8HotIapsZVO
wfivzipDFLpWGGczxAvXxGsk0YAOQxa1rYBauFMQ+gKgoS8X/68+zMA2gJOqpDXy
bzHlKlvTi+qrJb3SVsk8OtThYskvPoe9Cns4OWL/2/2C+WMGAV9wXsjfrogMR0BU
XUXOEzP5vDI6G46YkR/Qg/eiZ04M2INA46EiREwx0xTBQw4fglmYpzwCuS5opnkQ
xf5H6rrAlaPD4e7pNTZKcdNOestzP45/R9//Qx58fIEv/mnMcwTLfdb6CZZZMpuN
CajWmUfyc7bIeeWHOlVVAVfSVb0ZtP7GW29lqlIIsfKEktW/PWXUFewUmGTDY1lg
UfqS++CzDIeTyHRCL6w1Lk0mC9xXy9tiI8UagOY/ve0m94qXBUdUy3TRvDCqxS9E
FlINgt7T4TDw7W+5gMLsIQzEnx3iNgxKUg8KlTJ5UM2YGkotcQGrVhE0POqdDoTe
mIwbVTQgj8Pjnt0LWBIMY11hZU5K7aWmIF5uN6yrjqj4zK41CmYfBQBuiqidv1TV
O01356jswt8hvyTblf3WnZRnt8ZARP+Hcfpp+V0l+9UuxUhxC7yQpVEu+L9txgbs
pBCFNejGmNG4sWbImoMXMZcHLDltr+3KhVRTPqkLCuMZIZpUn+XxeWY+/kYb4XA6
Y0owP+q7iRR0XKSwJrnSF3J40DlYEBUv05NBSh3Hld1Uue36FYsddu0pGrZc+px+
LoLa41pq9ic+zrPTMFonsUKCWqxUhD03qe0uOYwTR0d3D6B++42MJsr6xb7pgC3S
3/NOnSeJ/AasaknBe/NUcYqRYdtnMLgO8Nxo1Tm8kZV/82w53Cg2bcVLCHOJ4WGs
HY/sjah6PbTYm6ktbGzZw512dNxpwh5CLAj5UC8cOgfpE39MS35EadSIbB8ehTVA
9fdt5Bwdc1CRvkNI62akWUJQjcmAe6LuI0k6OIP+aJ6QLJIP7SHKmwsAUP/HTIJx
BJxhGj2dOLCPT6+XCvS1yJoNbuc7Kth34WPoVmFHwsH3BrmdFplrbWqQIXEtxy1Z
BbZ9ijAcsAYeyPjCguXcwzZ1hGbm6VDxa/KSFSxgu1Dr7daUEEMcmK7IS5pLu+KA
s7sUmC3Pnito3/3vV0aws6bYgX9m/8/GUBGUinZPNjJLU9QRCCYM+9zHVG29ws7I
KrSPk8Yo9z2xUKaMZN1EVTWPT61Jj411A/DCkVbjQihGudwr8QzJad0cRgqp6ViM
H1gVqbf5FuuobkbFah/D4l2GYEgdpTlPWg527Eps5bHx0LI97q9pzV26GS2plIa9
67ixarDl3JYSrJkOyoIXrScTW1yNzzDbMekDLcUcX2+ndi5jLWhkQwK+ZsPE9F1P
/ItBa2IB3azlNleGaKCIG7s99Ly2kLgIoC08YSXz5nF1b+S96PWEcSukej9coxQH
GUtMo9WGB28bfYNol0zRCdD+J1jbJoU1eKlzOltD/6c/HEzwdZ1i5QNGNJQvTfFK
Mj4s9RK1VnxjbDQ7PgHYhw/JHdCljEuNEMKpnbKr6/s7WprGN17e1G/FZs6Eel76
soNUftXORc61+ceR8mjOsCVcH+qf4ZmdVK7KlmqjnIdcaSwqcwCKczotTOxU5XgB
L3s5SiizvCF3ECup/cSTDpzvfme2jJNjENwe8H/COChX4DWpVQGA9WF7xg11AHDf
oF5Ag8ZsePOMhy2Jv9W3DM4MNbnowrxSrp3RMAi9dQvqWgTQipVYj8hSzrAavBjf
8+ugZk8+qAHQ2k9xdyNKVeGS2izhJTqPtKPWl509qPauxHTfnG426kUIhHBilWcf
wLA6BMIhKzksSH3R/XvvgJXgqJHqwukNIrFo9pi9w+V6/9NtWWvFseOe2/e8p3dX
YZR1QiHj9datUD3+nFLW5EvNjA3mJjiJ0uFx7D9RTfb2/YDl0QuAhV8eO8bsk68M
GqX66qomeFXibNxd5S6pr892GuCGvLdtxED/ReT9zlgtvHuzCMyV8Pzd0EsbkQZL
xfnGK56ZLmIostxMSSNyfS0dt9ndepu6lu4Lz8cbs/7MMnAY8x1JKAtCj7lEBFVm
ab80JLkK+vm/JUt0sGqconeFQIITZWIxXfggOkHgrv+vXCJiwaYyy6+9rENNa6Gi
XAgfV9MUugD6ILhCw9BZuo9uDbQouAle9EhogWa9qkDMgeWRg3oO3ZtZybNnz+lD
0fNj+zrTTPDch6ylGwCBMnTCQHBDB7/fgz8JXO9E3hckhsqmNo2Urd3M4FFPm5Jm
KP87vLTjdMeDNQp97stT4K0hbpLXNfnxRcxntjXgOnoCBVGXKF5LNJ9WjS2E8YW0
vbjp42HSqpzhUcR1vNniRw3BaaAkznzkDHWa7v/4MHemN0Gv655+MmamduCJfxEQ
ugVy2Esqt2taISacq7ieN8jR1jwkJAJ1lKwMGmZt5jw5Kx0NlUuX/M4jWFqNPqL3
vd3AgqTdVnVeitymyijGwFTM8G3HsnYWPnQJFw0vUIHPQIRMVX3jdPlnggp9Cj35
FynxU/4KujTmCNl1zImUoOgt9dmbIue22C81SEACEvgIQ9/8CNdBCLpPvAAFoTmI
R/rH73zE9nS3TLrpMgrFPUQfUGCeP+iNJOTIqMHHY/zYWrZJeG59EqscSb1UtZaT
y8yZBWfPbiOHYaLRpTn10YkAXFZawqLrpSmxmkxLYw5wL+Kxzm2hT8Mwgc0p5hFv
y4SSZcL6v1wL/1BDDgCq8NoDHfc7/FubbcPpEGrpv/691aDtrhVYf2L2/ID1KMIJ
DUXFpuo1ZXq0j34ugf3kuLyYff1yAxA9d2nPnjlYKSYqo27QQSbjz02QrMGkyHLq
swcrSHwsxoGM8FtXyMHEVzov1OZ9q3Vm/kiXLnjHM5yR4tn56IUph47aV6xPQChD
tP9eGGc+deG8OyGVnLgFaxEtPd75WK/o7F2IrbYUQ4HwEPKBuINcDe2P/dd8tMSg
NeLvUpIV32YHQKPsR5ExI3bezCFWs0rnAC+/P+psmm9DWVDxTtR2o2Yha0kB2J8f
gDdEiWLc7JfAqnAUhpvfIp3kd1721SLdV/5KAFBanoDTAi8TYGKpE4zB2vRXH9EL
hlGtAdxH2X9sC21KC4HJNGZSxXjUMJhub3vUjhb3yurJCIyMsU9ZolzCNG7Z+FYF
hPins8Ig39Uw2qVzdbFaXRzyKvYLmZwMS8cFdfrNsp+Fs1O0IlSJzi0BfeGDXxn8
gA2Hrs10h62OlyuCvjoHCGGDIzeo+pEPx12UHYEJ6eTGhFLbsMnOsyHEkLAMfbMQ
7yzLRKvOz3Tn9wsGQT4BqLj8pDWcBsfmWRRaAxOTAn3btD+nZNOjWNz3L1rkLU0M
wbDFMfYGRBTQUzway/D2rfBp8VXEqAYixqKLVkn/qb6u6X+z4WGFutwC9V9P7rJY
mhFy/R/4T+zv0DdgcDhbMytCSYXeqtJeJsWmu9JJlUPBf2DEjzu1DUFIlpWzwn7d
q4QmwHi2/hzPyntBMh4LIm5CWJ34VRLxPTFCAk37KYGSbv6zscQFvK9weQBDZchf
pkjR6qB/zgdJjh9iGlNf1nXkPld6FA2X1iNhYYeKnp1vwVqfEG9dTFHvOX/4KYz1
ksDEngC+Tg2KjoHMjCQY54xXo2lKIqLuHKpEb+GZ56rtQHQmYE4YfryWj5MYhbFG
zKKz2Abso42SEpD1pu1Tod31iAQyBnrbg8kNRxwG+0cM+rlOT8tKIJ2gh0uFG7j0
cAV+K+ar5P5aravHgd1WZDkKNohZDePrLwWESA/jyVuWaJvlkohTFDZJcA2iMhQh
FIASrDDmnkx29R48vAGdtRIQYd4XTsDCJO0q/JiqqJBtGF9S+0cHYxhdTOg9K5OW
IJrRtIBkXrqodKIvNFqaNPn32rNYBGW304MebEdJDADRar4YfXy/3uLuFu/Vz99P
fQelm9P0ONqcTULqdp6+AEVSzMw7jV2MjKNy+jYfOCLRKjsILLPlbVf2/NyTkJ/5
j8qlwU4lz1AccHxAzoaVfDePQeRRQxjeQuosR/B2hcvjJwwkWKuWe7jj0RRYBsVw
T8+Rvz5QUsxrZXv2fGYMwaSbLqJPy96qYTsTPncNmOeHfYe+MgbRKfPDTKdVIrwl
i+C2BkcomJVP68nep16z5gSixB7L7f8jv8MFH//zMm4acSa2X+Z+t7VeOOhZJoOf
aAFEU2OqAaWh9a5Fnn7ELhv9pKEqx4UXg9aZ7oMhwYhGcL1ZNrbUnmZn3UcBmUIE
74TtZdlg3IxveHS/41xQNpSFx/ogjAeb3vK8SHiOsyBe0ltXoXtoCitwpeb9uZh1
G7Ja667GVxDtUKktY8O0YpKnKxGCn6mfAr3NsalNojp72pX1QMBh44uXpQvV0a3w
12V0KOtWvh4ElYLhFJq/pJxI1xu8J7T2yigUdlthc8lldwsE7V315xb/EP09Qsv4
OGj1YXiVZtjSXQTtyIWExAKoylDHKZmcAwG7FB23wvCqMsgKWE1lFbKifE8H4nyx
Wnyt+IMgJZA8lzsJ2rRJ/MkZmBiAVxRbAOs+g7FIQU4sdYG97GdNkdiloJg8RQR0
hIxPIPByz7dhK7W2CHf0kw2rn9UfK64yUJzGS9NmGShVrmj+YCgp0uOvSc1n4hK5
vRlY8S0FCutr8jLzCJ2XEOAyiMNwGEsg9srzvtLYI/MnyvrQ6k3MHRzxSmlmrQe9
vHXsJUAyoS2ljW8P5HmajnZoQwEdopHwvCwExHlLy8EwHscVZ71OLHGegzsFz+39
Lc5kUBjkhb0GXCB/2WawwTckduzHjmw+leZil8qMo9a3zp9UQbLBO0qhnPspI1cN
pWk1DsD6ZYg/uJIlWqvIQ/5jlCdOsiyd8beIygQEuihqBloVEo1GKTqeBv+7QgnK
jcutfJWPvYla488BgrRQjvwqe/XUKlv7+vhm35OY+HCzhRLWS4pin2vmlXilKVA7
Kisa5jtjeJhnTW+uRLOCsW6gqUicyA94vtPyM10ElCIWgL5IWnAzNXazhGwj4jsu
cLHBrPNg+4Aa2xPgvpZys9buvtuCsfQbN8m76AUcYp3Ku3o2HCppAiubx+YWiVdc
XBDveTiIXKyCpHdX3jeibj7KBgbzCtGvVmBLmCtp8ZDXif3/AKxxSzWfXBm8ZLCB
JCMf5lmVzEKMOzdJGLNqDWPDMbu5Ke2djrXCaO5kLCq6ehOl4HTlZ6u8ehCwKwU7
NTzm7kQIn/rr7oBMWKh3SnBayyY9HCApBWGT0Ynj3Ryw3wCziISaF9o3PxWNBqhv
D/u97mwgVFBicKRr2bL2VxJjWgrIilmvlpVd1t69B4jvftuozTcRH8r9PWL3xMip
LbQb0dWSLuEqwq5vDL0xiiMjmTgkdUKv1MVMrBXtfCXWkrTcXZx6IslipOcZIDWG
wvjyNZgI6eWK1pYEK82lntSdgQkNYerD/OurG81h7Q1kbtav/L2cNQvZcq9YkYwu
Znbaggm6OGUc0rE16iOEA3qBg4jfkuE3EwuOBi83DZJ4tF1KGSOiGmSazVkAE6xw
rzg2tyLSnefVXBoKRyF5vNGeKF3N4Gkzu92CnatwXl4X9eWrlmHfZ91k2ofTWU/q
PMva/sCSAiRMqNdycodypWp3NILDM0ehXlDn13gyF4VDfAKYWAcJP3eHebaJT1Pa
SRzEDI9/12QKjyX67ORaAEU6Y8LyiwR4HDoAiq9hHRdOJochK+65qXGNMiSiD27J
2QPl9okOcuuSQ76vN0TC0sDeP46KSqBeSQ0CveMmzbvIoJ4S6StmP1XSPL+roM5Y
GLwMON/OV/ATn6RYuPJaYRR6Eah3q5ABYvp2Em6c5OJSnLSgts8N1d/A5Y3X3bUx
9YxsGs45RM2kzmwk0XI82J0wPMv+lt5EhuUitu8ePtaEuRTs2OgTxhAC5Ba5Q+/r
p3CnhtGlpIcr+HdTKGYhw3dwhFwZ1XjzNUHozSwc9Zzjlia1RxxZKD7KGyqYyK+C
WG89bjyui6HsQ5nipPrOGDcNHhgdPkaMGpABViBwhzdQOjJJsHS7/JuApQ6GK3q5
+JQi820L6Ax5G17AjhRilej+ZRjlPrus2U940bN32XRSk0IKqPG3TZ24LpHAmsqS
Q4XSDoj9dW9O8puMkLtxgihJJ9o0lQW99SdL7Lkk711P3XYMJHnL4OeGF/5nkgaJ
/bv9GVaFTtMcbQYnNLbHeJAfI3BotzhbTyHUQ2MBtnjCAIAFy0qTx4hKOvxzdAM8
+Dj10UUmjL+HUiGUep23KJy+XB8gAvn7Hpbhukl3CjkWSqYLhs1hg1SkpvkjIvHA
dmvU9bwnm/rVvNX9T6eMXy0HjlZxp1KMM9ERdFYgxvJ4reMX8Rsr0HN/utLd1zyK
O47fmbn1xbB06H3qPz9BiK3J8emsv6ZmKNyPlorVvn0kQsGtv2xLOFI2v/hwcYNo
hweBQwMfDeZrNXE/C3MFOMvhb8DmmVMfG2WBT1TZUKfhyKSB0JHZmoTz77mco2gb
cT6yjoYcAT2/mHgqm3x49V2mYJZ8bBH9A7l1y8A4ooKZ42TdPkvSIShxTlvZ31St
ltDsP9A8aXzv6RbbNNcOwY7wW9JMRDkH20qxXR3tm0JZFx0RCNsZxmkYKUbVSp5T
/yG2JdyPyrnDN9c/Fw14kKfwvR5DN6ZOJSInY31u7tI3HPoe3R4OORgnuIHnUmGr
7Wd+xgy8HPK57eq8GtQi1TrC/bMLenwouNJ4yapomxTZIKkqHjV1K800yT+3oTG7
cD2x2Kg/I1PgGSfM/E5cxMvLPuRAQJEfPptJLQLa6sHFAGUuajJTbkxmTcVTibxu
2AlrszAZs/VgJ4ioRyuGvQhjHp95bFiqBcg/6OyVQ0hjjvC/CIRUNIFa9f3T3twb
wkxtLJvNj7Av6h2K7sTrNykURk6nqRnzc2Mvosm0bnvNeN5OIjcrNPGdlgIeMPcA
E469ZDmsER8WQ0/78SR2PwQCQquqwZBNX7finWnaO4yl8ESq9obnGHsb2b/H/03/
MZnc1GfV2FI+i6Eg7eDH+DbGacjuMzGHj1LZxbfTJLowzX7Cusx8ylvdoUSnCanP
YoCEh5fZbKo9cY+HNgSajXIV04WTYxVjSbYZTpj7ACA2mLjIB6+Ca0wF+Y2FbqBv
vIfXvVVTmdOLzFlD8TJRmKV3wMgAV8h1WeEsUqjWHlhsSLlebj9cxuZe1iicgZ1w
ZweEJGqoP81UlFh2W1zGKy450CubfJpyP/wQ5+BB0vA3erxBxaC7yEwTtulIEWMA
50RcW22TMrrS2Q3b1IOnePeeWYaWqiFw33+Vq1OMBSyiwIozY/koB9T4NqS9IlJF
MQuxeK24/HffehfY2Tkt5adNr0PFd1tY4l8CbBmmavx965LaEiKEqppzwN/hDu+O
upUFOkdoOXS+U4U3Rw6oHVBiUBuZfU7SKqcKadYlFD3SD0jQ35QJNxNbMK7dO0Mr
4YMnjlQZOhUfIsSD3meIy8+IR6iQCwNyoT9raQvXE6SrOI4DPZie0AQ+grOVbNGB
3+kuFd+iE609vXO/h9M3mMIl2SURIYiQpeFhs1Z4rD8KvTKAIEeH4MmpEzriF+/U
5rXpyAqsf6IHp9oW39K2vqu68iMmHzDX0xNR7NZYLF7h/r5GpyW3mz9PSu/cjeRx
LnMiy1ThgwvbWCAwrwX35sT7P+PpYEPlEdIOFg4vzrA+ucc0+QDGwmyy/AZA968B
DJ3r+Rbv3UmAQAxDhjPGTQhtfafa/vh9k0A/mWBxU2xOA01i+bHBYgDJSUIOcJy9
C6MLwdOxUOhdZFkLvVURTP3TLf7ezU2byrIGtxcFt3IAGd7LUHWkz08cuiaE8sjn
vF3YxjcQqUSNhm09HmxCsqTjndeZcnH3vdnZMo7ls8vO7DGblaPr6V4Meg8VIzzL
sEIFWKKwZ8LgqkFhCUYleV0dgcqH8oatJbEqSVR6EaxYty3eq9BO4SH2dfQv/JK4
UZQ+zG9m2L1O5oVfid6sBwQh19n01tt59aP7ATMvUJV0MuhzQeM0Dc6BSo1Cpn2w
2Qv1ag3e3VEECA3sH+3UwCD7nDB+8C0lFgabyuoTzNVi2pox8UFohUby9S4fttku
gaE74xNecK9KVwu9QW+fJlSgB06jj9UyIOKeHHQyw2yQQcQY8igxS6feYlRQsXZi
eqr8LctMSsfq8rUdVpQ0Wxm/TSQ2r8FJD8yab6NO2A7hj4+mWMZducu58FOPL2ua
36gAvUKEAr+MCIYHV9s3QE8xrA3EHhDKv8gi6BDqnbQieMQG31jMjSgi1MhDd7dj
n2a9W6gPga6TNm3ZHWXn0wasSwaUYVvYR8052xceA6S5YPCRY/vmGtDWQL8GeSCd
/HNxmD+zPB5ZEoQTbYVPFVmo+9HxVspV+1+AtVk322lTlNg7huHPmx/5aLIV19+y
cTj299mULkbR47LMqysD6cLR8SvMmdCRcPiw+N0xmND8RqCdr4m3hae2C9vbkh8s
Uz7L4amOs0NNnASH9yj7Epw3IU6vI7aKnqYV/8k1UIAA5TRZ8QXxRsKfi6s7iw1C
M6jXlaQDw1wkDDiKBvnYqXXE1nlGv2IfzcITuj3QERaccWmX5vjHaSo4mT6d3PKg
29Nd1Po/4CIo5Ev1jHt6TU4v1pBizZMAHcg9O+Z2wTRo2YCYEbb11ox3YlTPgMcs
wrVMu42ZCPjIPDE/b/n2eqrw6IC+5yFkNTXlTVI8zqXnJCKfeOwtY7EwCabevkoB
J+xqV9lvdOXr5MMGwQhfgl8CRrT782pDnPJmNBZKCB/fq0u9Y9OYeYXK835QJ3IY
DlQSr6ccwxdfoSucaBflsvaIEI56QLqhxSjZGp76TyGE+8OtrBpSND4Yk3BF4qf5
tRDasYfv4LO0v7MtfPTdteY1gMgAHwuITkc6IyimxP5lPw7BjD5hmhQ6RYHI5Ou8
g8lSVWQ+1O/wLGABIxgZpmHEx6Zg7oh/54fvBLKXnt4ZgPoWpFH1bgK3Y68h0/ir
key9GwqvCSICWsxCsR7PiQRH0dzDqpMDRSuWSBAjML1GFR73bQsFJnymFDN89Otu
fi9l4t/fR+ikrGzTp+T0ppJZcXE+nKfIhZk9QiEF+IoaEG66UUbpcTi44DfEue5E
QFC2HyPnV8TjrvX+nUA0PGlLthVjDaSVe14FYBxo9cm71uK0kSzjJzA7l2FBXQie
AgeeFmAZczZa7rN0DQEHIYrDrDdC1kqS5xuhBPISvHoU3mnATNVJQgg9QDEsvSUw
aXc1PiTPx0O6GrAtX+zcWBhb+yy38YoQNE+g60MzBBqBokqQ91dSnXglF5ohvsPG
oi/y5NKXNHiVgU6jiyrH+RxxhBs2Kgj74eWfEHEKWBSJTtlcKPTuRzYSpUnhpvZo
U7bOiW8haCLuWBdVCZ2T0Akn22CwWd4JaroU8A3hU4XLonnGEy/mfzSOEQeK/1ZQ
2VAk1tybSm6n7nSSZlliRDEXZh4eJjtjHo81/1EA6LcF30VcNVs0R5s1BdjqdlHt
Y5I2mLVy294nUwnZGeS09rCWfrvFQqLD7jifWQStKx45VULe4wYj4/69MXFIpWUy
dwfbqASnrMA9i2ksioWz4abUU3fpm+KNhXarUznP1G6hGrgSz41EzS72sPkM4hHm
ffHf2FqJCpSKAceJqo68nr4YF0hTOJk0Y0lKA0isnd/5sUqQEU8a94IAa5WIlEId
Ayh4HXNT/hoyR7HIMCcopb4dSZe3yn2FDPZGC64aK6sAzYJqghpmn5nVrK2mVrJf
HED5u92I/1ZaGJrtTnGMKDJxqhvdAsNKdd03feT+gR6DqJC+Gwuwwv4pC0ybFLWx
uO9zwJCw7d0JKgaSUcA0QBKwaczraiy2tHM70vtKSAw4ZA3DSE30gLnxPmI0TBtm
R/E8ULJaETQgz5T+wZ7EMefMqOyUMpskaLESx1qltC7Xs5a/AqSkhKlI12skidPd
JnLOKRsMt7LcrGg0T3Vbylg07ar79Y4Bo3UYLxptaiGErUEa6WhElfTx3xjjKCXt
vGf8zn4CrU+a1Hz2PYQXm2yxgWSNc/ixH2hmjFG7+LAl3T/mz2M72Ijz8sPynxtC
8x/ifW3n5l3355dElBJ9YUirq8Ce6z+nihaysqtkzg/+gAK1mLChlZ0iOQmv5aTN
Inutqq1Shq4wYS2uB7IHOqDNU5pvFZM8vXgEwPY8bgpaHwjci/y/zkkjbzZtX+x4
R3/zrKoLATvUKgznGmh3O/jz3Fk0doafKyhkui47GnIFngVg8/rdaCJnZAZ/ySWh
EjWCTjHEMHQ4btpq++UKCYVGMyOJCuJaHd99dYv5UUYEUTnxcuAFXYIHGCLBDLzc
wr5FKhpPkJgivW6OnomQQJD8F7kP/Wyjrbq/pG3bf4ViT4FgfuviK1UGGFLl3Y8w
v1i5hOg2zEUsLrbjwxHn3YhGNiISiwdX74EDsrku3rvf78Zz1XFwEtRoQG/GO4C5
jTVLq5IcL3rzUOTDY4j+w28SfvBBCyCmFTxXdc1v2NYVyenGNASLPL/G8WYdr9sG
tN56vid0VwFWIs+Bbp51SLS3mSURoudydoPtTrbhAI39VmrrxcIReiBY1ijJsZPp
BreRDY0PCmPXWTRIJD5tghAoL/gWI9IB8pZyQCpvJmdYuaoJF+Wd0Q/z5XKxdi8h
75zPuJiq83Gu93lLsgA66UKx772X5gJuZSnbjk7DDhtyUOv5oYkJ09938hgDcPcg
ShdaR26BufJ9c6sp//lARXqLO67mDvvV1Akhju3gTcaFqqc/xyyQmFi6uDZIWKun
yroyF2EhunDabicKkc3Ddp2wrR9SjYovqApu/qi6BlY5bLJ4jIW/hPmp/GRFu7dL
YogUr91gO0QcDeqlEpYYoiUpEeNbHjUFoKcIzTJoHovyvPO59Ptq40iaHHaMitnD
6RkvnSRqFMmH9gIQKj93Mj4I45CwE+7eutbMaYOfLtcp7HS28Pd8aY5omT2YUnHM
mJv9dJaMLMzbuFPDqU8Hz1diYc2hbgzsVDXdindIzCzSvvGpVnOsEbgGR7IikY5w
smUzJlT7dKvpxkTz55s9ismFFgJAu5WLITSFtPXAkzybbtDJCBAKWriC3sC0kbHN
Yydrv8rDaZUcA4zceBFNzIzRqdkyITtNIlbnvd5W5zdk+hGZQuPJD3PCkUpVtlth
TLAGzDHQk5Wd+UTLpsSsIEL622gsrbhoAftE+gutpDWd7hJPktiaCCzkymAMLNmi
jkMrGawnLU6RtSHR5VnhLGmKCmNk/8Om0RBystGC5N2Bnq3mxs/gudc+mUdboheR
4VVS48K7wtLDMefkXAAhxUplbF/OCEteezRpVyNFRpix4Wah1Y0jt5lYdBdyK/Dd
mTnrYs3z7jbZqf6rh4gbdswCa9LrQm9EF6bpghgRHqtILnWbBKjIsSCO4mhMzGwS
t9q/Vh17Na4Br0lBYg0IaJPzlUAixpprzw94QOJ53Rx9DG8vaBB/IxPMA4/FFVjX
haeW1zOc8TjeHeHA7EB+auAdiZVoKhqoDMeG0MwLZMmNyKEVe6wsy5iQBAumSthD
Ig7q95brC5eySwhjhZvQGDrYvjzyBn5SwT4Xp4VcR2H4p0azLX0rwCB2OUAUzaNv
sR/X1fSGi1/C0h7bnNxvMymLCDfq/pbN2aSne7V9KucXPGJftSjGbkXSfXI931/L
Fd2uA5LSzb160C4gnAm+0eHmJ/uIjC/BSAtE4DuJ/YgodAd1gJhqoKpvIidQvVUv
WviQmGITXKKuOCuWFxyygOJBdSlkZsQc4c0Ek8R+834K/VfhIgaTGm3T73lNPmQt
uh62Yeu4ez3M1wNLbwt/oawjJQyJqLkbajS7aEVpLk6HjG7qvriAlUcb7apPFnzl
dEoS9cFC8X70vMFOi0KKtV/9Ozvgoqq1lAeVpG34n+r81IAHlb450SbAjspsoTlu
EAiaYkGXjK84aQnqLYfkeTxIuOrw2viq8yOP7DAvwefYQKJhiNGmLLoUGzEIF+FR
ggKWhMyB2uGbhXFs7qIAHMoV+EAgDI8WVTh1P22jddc0lPuMBdacD5E26PckWDxE
UUwQqVmy5txVIXw6RMD2PIKMER+qLg5W6IyGVyi9IlO3VX/iJv1IlmRwtsb4Wo0F
QgJ3nD0onhhstLaCIL3Cz7xo45ljbp8mvJBBK7g7ZS+9CaesWzTQAvHjExQiiOsx
8mTvHp2b1DykLkoWDvzy2r5ClJa/ZLJQNUBmTHMWPB1HZcBZMrPm2U96QcNZjnE/
A4oC8J8vKtzLd9l6de947RJuQxhZwNqmC8Rbwmms94g3anpH32UO7fv/UMuccWff
3sMzK+F0icpHCbvQeUXlvdhI4mxCPtyTXVhQnjb7wBckG/mr3yxysybyXse9a0FX
xk3agOW8JYXjJRFMG8WhvhF7shT8EXxaSSG2XYCUc95+crfs47r+WqUPwvw+lyS6
HVuklZP4RXi1IDQqNPQhPUsZv2ez7nqLX1UZVuBTcu2BbPJQUOrfLIKbaasFjb/j
MTbliV2Yu/DX0blZAlPFbYsOToVCq1yqmX8qVMfkq1I1HqJu/xPwz9MHtQvIPvGe
zkT1uu9zvIOaL/1ceD6xQgqqr3JNQ35vgZKv9hCpzJHl10HsHxWSAkKNb/WJ5ueI
ZngRQl5PcYRulx1rEj9RJJ/cF3C/mMVELXCHVauSW+G3b4Due6hBlAK84f8mQLU9
ZLZgZIr7Wwp9vWa/ovpbbFKoEUBRNn2pd1LL5gbIZ/IVuKzpUBzIMBN7WR+hJDR/
k9oprweLs6iF+OQirf4vpXSNxeCYDA7BXb1KXLNQsQmjf7ou+fZ1ZClJjbfNjmTY
6ZcJMb94OnlBuz9hKuICIUE74on86AYaWlWkQOHdkmdltIHY+3YOhiS0k3KCaEpZ
G6c3JR95PLGdI6BTcyYmZMPm9atbMtzvNfCSYcA9VEsz/lrpv+9LwqiLRZbfxWEx
6b+vQMYlw3V6bIOmDD3wUcK1H+fcJ9jB6hQhywpJyfJ5As2SjcDpeKGrHk5agSVj
Ye6D/iB1U+fJbzPp3QzF2IT63rTkO6T+4zxosOfaOlEIxmSMki4FRtI3rfy41MoJ
JDJTfottVOX05A5+Y5fa4P+7gOJisyURWh5Q5f50L9HWSZCMOO9AFYx4Vk1RJhfF
peH6zP4eKYTFUTzLcDcH0fQT9i+34KTzH0e6BaahAJEsGJzpRqyuH/9cDcxo4kKp
/AQD3N54myOG/xHfKLFAR0i1N1XZd7G6Vpv7OQKXfwwQTCZtf8mMq7eTjXq5UDIm
q+FJYMQfd83jEUH2PEFqTr+3K1F4Rlv9pxCPlsxqfbWEnY1HJ5TYMDlG+zYU9w6N
WPkNDSloCj2klLuUX9SBP4PZoFfNU8gIopDeCWidEsiYThN6UKbBhqR+s0sNjlMu
AZAySPsT060wYlKNsGzePN5eqiuryJozJyjWZVAOlwx1M3/77Gmk+bo8wFEbIZX3
M9LsXbimz0qQQblrp/RpVJNJiZE+21ICwTAw7jtxBnlWeejPUKCtITY2Qsa8VLQb
VQWzpQ83QHNtDprOLe44rXNiJFHczJX5BS7IGflkLTTjfovUiFcP1Z/zuA7j6NgW
bw8hx7Oa5m5igprvIo2PgTY7cDFqS6PR1FaYCT7Vx0yGZq269sEBdRUPgdYxla5q
WyKH1yn2F5+VfkQqf+fgHrRv9SudduIKZj4UeesGy4cLfWK0/4L68VzRwcQ81TnP
p4lut3G9tsCKWeuK++RLWfmavMNVEj8H+iNhkipIV1lxC5vwcgId/UOg9kJumDDw
v1mvV/FFsohlazBTgPN8a2610DbCSZZeLZNkz6xgFATuRFLr68yRoe/7ZgmYRkvt
RzYRUp9WsNRa6HnQwlw5lduZhL73j1j+rmurxfWMWSQvswhdRTieEQ2mMmsq0VGm
ukTtQUGX5XxyMWn5uuxGtTy01TrOsQXP5zcBmEWIbyv6DQLbP+uu8vkoaTadsLZE
r1rSAN34mFtij2R2vYONqIwncY7rqdxqNVrNgbKvyLK6tMizKndgBudJqGFIxkTD
97xeB9UN7gEmsDwh6UcXhPmY1Su+546AkBEi40wLSPtToFO5Ipm0J4GLCXlTuHHT
jPYrc4EbyyKVUbApQL8WAyfU0nEUu/uugy/JM73xbYMlheMW7QSQI+gj74od1KkI
R97/n1GIfRKMkYNyPIsQgubf31fvVrOSpZvN04JsG9/Lof2LEkNAoBoojSxEzoq+
WaxbdZcq1EQxhQaXThp5Hfhf1zSfJBrwlBnzMSBpCYdIzvY71KPry4XtxaML7lWL
iVu+Kn/dNCv68he9E6WMx2Ayz7UHakJ43qMoDrBY01RSbRc5xX86rtLXwdEmV1bN
+hy0pv6QfXB9bnTXGaFdnGjFuHAKo2Z02Z29wqWxPQ06J3hMMkAHAgCwcvkg7+Ev
bNXAAjyYuY4BCWWEFYodtrQwVbzJRbJJAgzkCR/KpDPHc+pbEdWSULO6AmOe7E0z
6fcwhzcnzckN17uvlas/FlX83MzrIypJF7cp0q8mxf1ojmLqLOeQQNnpYPXSlWIq
n5fw1M1rK2QjUyHCyuUFaNSQbn4wHWs4TgUI4hI1TvUDo43piR6ah/VuISzzZIdQ
e+tiT4DWLgUhOrK6Xfgi/3UmO0hNeLBSKp40rKDz0mAoFlhc1UDva0nV6TvXRpxp
d9Pl+p7zx/HLJQ58XbBTmMGIUR5prHPa4BKnm3/UAOMPkX4iBdufEgy8naRbTN8I
f49SnHDRcn6dQ8HVMmf/aFpN3orQ9VZmybEhDa2kRRhI9Qb76rQrzmUzuZyg5iAi
KZVU/9EQaHsgl0y8FK4z0rz/2eNMrXCaFycqfvpE/WpV3YZgInXSjY9V4q7ez4gW
NPbytlv+9tGSRMTQ/5urC/JhLWR8cxi33PkcREsgpM+ONYBjbi/cSrL6/GHubNg+
m0RX/UpP0bC+b2IvWTRUUpmIoKh/6/KVOdcKxnch468/HVCvIN7oLZKoeCmoPNzw
ItMFg8UVW3nmjRWUouI0qZz9Pr0NkotH3c70T1QfCsBuHDm2tczU2WGEibVQM7im
4dux1EfVo5m+NhBlUgt7UM9QWGqexu+e2EqEJJJiF/ob+3Wgdw1QXF2GEW+6+UTr
wyQd3/oQtxH1QZqzzJjehNLzw8N5BcIueUPszUS9HjeMCHts9Yt7/i1LXefx+VwM
bT+EbfO+oU+Vvk7oNXlsTYtZh0wIDDZSExp8XdU5xv2FwV3yve1cUeaHtVQFzhWM
tPJh+Okp6Q1P+qc2RSUlBMxXeacoxnSMJWF57GD2V7S2DZWUQLw/TmnVzZyy3mCB
BpqTbrO9mCZrzv3iGsu8EO9Q/qLS6Bq+EaUz+2uHVp/c8jeWweinmKdGBjO8cVC6
4NRqGW6hQQcZBb38CFl8Pb5jRKYaQknVoO1TvEefBJrbfvkRpJqLbatXzXyYKHDP
ahulEb41qfcrABeknOBGt3n4VoFeEkIfBMVET1Ne7F+kbvPrJJ2eyMOO/abZ0geE
KYMep9OcH6LvY9mRa7IsQnobnt7WKOhomwuXnoyoBRcAjAwyTSNg06WN/jwrvS2x
dMXloEDIBYuo/qYwc23T8x8iss+NJ370fWOjAiiRo+t1hzjz9ZJgrIQymlzZhdpZ
/qEquBn2+V4kA7/vw//PYWYhjnAYEfn4bxgAIpqztCnHBZ0D+p4/0SF76S4rRval
ZI/G1j5LWVFw1T/8G8Y5EoZegy6Oh8qxR0RbDLMDbsYEN07Fr29IWwd2lKRxV1fo
a3HhJ7Ae1SGRH8DCXQSi4iF5PfK84YyjdjSivyqB6EXx7EseZh3R5lyNpbhrB6gS
loA9bAt9dir1/5trYDIFXxX9gLQlo0MQvf5C4uXONHxe8N3MXpZW2NtvUzFbFjcS
R6/tYesb0Ag5leDI1u0ZJ6bpxlS24ypKEG3/caILv2uDbTuuPnpTGi383rwsF0hN
Bu6uED1aAQ/mImOkuAw/sQTVGFrvgwM4WVCs1S8ZyBLxzjfnlrfJ9lWxJp1/PKOc
g0n9CTLGTsT9Rct4g4c2VToALYPPxMh3/4iElvewOusc7Jtp4/95lCNRLzODPUu7
/pCT3zLkE7u/D6rL6qGlvZ2/kOulYvJiIqR3HDr6YOMzpygInyE17l8/xRh1CMyz
4/F4eJdLHOj3YGM/gNRHI1HmvgfKKbBYIrECg7s4Rq8K6zX5Y7P43HO9Ubpg16r/
Fpd5AiYxICaCa2fEPmKv9sykyTD3vtbP3uH5mJoVt9wi3lq8dTzG7eC2YhsqwlKa
4J3OirxL9800IdkmfQbLH4Ow7YOMLDBad2WZex7PU7h4iDVKeuT29fTA4pDYaVzN
tqVO6nQN8ZqwCwwgzemBRxpoeBbX1TJDj6YMldYOOzqHYUq+vl8PU4inAq9NMOZc
itLtyvTU2qIFH60Gsfvvc+oNLWss9ZvNZQSk7u3G9tKWws+daI9ggXloO79SY9mn
pGOEAuLbnoVrvfaayRd0WvyKS8kDIm+Wh2O3fscl1eZzkRni40GPjj1mzSMuew2l
1GzwX5dBiZRRN4dHozzdGkXKdqJ+41VlbOft2f9hvLuZOfcyi7dBAAdR7LPs2bev
ZMORaljx9OG21mRTBd7XxNnTnCHJyKPyMU9kY1Wb9rBLpz1n+B2cGZRa6uB09VXA
n+sMtNMAjEYmQ/RJbHOHzfGCixx1FSSRsDscXH3IjhdcIIQ2vhIPFM3eqs3EEmg/
i7gAXU35vwPgAO2bVeMVhqyhZjGIIxBAdmCEBBEZqdcJ7pBzoVOOVD4xMAw6FRpe
G0bVMpH70iMd67Iw64oGobxixi/Hbd1SjoF/zp+oMJxILkVZ7TuGCcXpt6WNn2Gs
bQzUZuhmzfKAwZZxtl585GeGcmSoPpbshX9B9WRTknEA1BgeRMP/dng+r8rKRSty
Tyjn+s1W3x0nbcb6qqEBJ8LKp86z2IChnKJjRRyX+mkcxPeQDLgQXu2tihgm1KpD
h00qgXmogsjTweTxmrUIWm0iGUeez34bH9QtkrKPu0BaPvd6V8HbhJtKrMY2jm8a
7rNHTW/YBYs2wdqsM3+lhp6kP/hWbjkcTMhPHPpLUVtIJN8v4zqAn6+leSMr71V4
VvOd19pypPHxrV59GoanafdDmss4iHEk2PeFUukiKpZLB0u2ImA8yRrXjlydZs7i
w1Q+zD4cs+1FyDef0zSKJxC9+6JBiCA2u2R7luef/rj24yTWK0DCMA2aTjw2XCRN
JXs8+ioubibw4On92YnMtfaklhy9QiY+S2tCpactHcLn4iej0jqPQkDRwIeo5V+J
hvc+eVSGVufgptlC0pomWiVV3NRrVanDYB8YzmPOOqfgyHGFl1ZXyL9jxVO7XdkO
L2hgze3NcsG++YJIMD8sW+WyS54NklDsOwjqbMsXrtmEuEF8tAbOmrw/kfT2y5IU
uwHyQPmkqwW9oW4Bbf0qSxNf+jwFpUGxE91CwqzxyXKV1FdWQ7BMOedDG5dXZXFk
SwJplVVwyOHecpruVw9c21KtcvAYyqv0v/ZF6BBPgCmqmuHpMBiKxvjbukZOLQo/
wbHwhytUwO6thu7KowpGpK74LX7f5N/qU+M8YoLUhpYv266VqsVelhixy9KnDJvk
ZJFqUQo1Ux6FeLtw/Kw2l024WLXczSt+2W5pgWupu+84jd73YTtjnda3Qhj43eaT
mdkkLam4va8YB4ycC7+5ZNVIKLKz+rUJItACmBkR4/QJELOiyboepS2DRtrs3VpY
5wVljSV5LmYLUBCNcMRJ5Sbbdehx1Fun3+YFXJo5XQC6OozHKqZHx4INHuswg1Mo
6AotCs4gI29QcKRiJt15acywEAohXZMNDlp8wKGU7cFcJqQkxdmbpneUT5YdvdNR
khDO1tn8KXgO/3+Dy8nL+pWxlxqYFGoY5wfrT0fMS+43q7MhktyXnbUDMNJmTm4f
iY0BkVZvOv3syc1bGgzP22/HM6VnzVqrjZzoa0O943grKR22ZLp3mDTm9h8mMlfQ
DFPj52Bfiykrc0jEd7exlzNmSG2RdqCpehDMweE27NgXvlJhqeUH4EnU+0r+KsMM
5c/PNYGMwNws9XxxH/gaqxQ/sHHR4yIgG7dECTK8CcuhAgxdvv/oWZGb75cMjA4c
qlunJSvBh2dev/OC8r/j9XSz3Eh8TuVWP339rS2CPY5duyBGPjgJUz07WBcxU3nP
5CKHXU4ZCyvRc8nGAPBSF00VRS1FrNC2DxmDzZYDbseO24+QO0ZDXjVUL0Zwb0pl
6m+MKyTVn4PL51dIMd/n3erW7xBN+OWJlV3JUdwZf56fAhJjlhBIica7+g6Xdqeh
pGGj7StV2RQb6iIx/U3M+beLsmi7oitxtSCgJZ11tE4fvR7qqwiJCG+h/5C0zmff
k3mDACtkU/0/MYiqmpFwUewjxrVbd6BEo1jfY5EewDLl2yXREI+8JSjhA6Z68uBh
7zPAMYu0R1xhkuMyxhe+4qFujAEzV6oYa82Es/+v3YxvyrCtPFLWpEB0XgGFuUWO
zcpAu+KP+ef/sQOLSKK46Wz4VfMf2Kxwo19aouUomNLqnre0Y2opBlfzplGFUHlG
D35aq8wqR+H1x9Da1tion0yrix/lkVowFjlLgqsZZ4WP/N37Wsy2sgmYYgChUu8G
9jE3NidyXYYzbLhQ9btExflzMAUUAt9dLM7oa0pBbIoW0MqkgXSlFHYRfpcF2yOa
pKXJUvgNnj4O5FhxtV13N059afEGbqwI2hIQRs6LaBnB5OIPN71tAoDp9HpahoHO
4/gE26NbKz3duj49DFJhkuhgB7l650AcbGK29FXyujMsVrVcV6ox73wBI3LtUOfE
8f3OpfGpTSM+WLe0jm3C0rSHKSxdakZWRVxHTUdGATvOnGlZCmoLZQcPqHN7LxqF
5pC4kp1Lf2nlUSujx7vgGUNR41TPcU0V9/Dx+yOsv2twESYJ/PJrBDdDtyAnBKLa
a37DPi4Cp9knCPwk0HiptUd6sm8EtFycxUPSLvRa/bfGIHCkeZuJVpzA9w3LIQsn
T9y8u9BHVIFX43kLfziLdHGvXspXh9GXWi0ayK2Kv5iT4bgwIlr1QWzcFl9jZNmd
1eMmCTWOy7JATJU7zW1AVC8LWpxXGLfbnyMRf5P/g1ON3BGksKZXShKaPhc9dpyH
HUZGj34hTXYodqTEQxGnp5H84U5jnSsPYsXoGhhAjmRtEgCSBMpBjWRLvBJIK/dT
WPinDwsXV02iUFYKNlDXBnjv9uI46HXBpGxhjX19UmT66LAv0cgH1EqT90E4w6w6
+haXonvncHphPUG9sA635TZhuTBEZXHtOoR6vYmRM74DCgL1FpkmoY+Cph+xWHVk
1WAlHJ0aHJcAWmly2pxKYT3xRKI8OHUfh1h+fAg40MFpXVPlHm2k2pxlrkfSSR5p
/eHNEwrCxSe+Uw+FEM6mhCMP3pVK+GfAC3TOVfzwtmKoIlZX7EckIpM0955CSteS
ufRhKRcjtAmUwCMbnoY2/zKNv9nDOBR85f87NS8mfIS/COyKdbUWYWOKPCpecHgR
A1IpxigZpgboe3/3neI+pYlBgxfHAwhB5zuraK2wEJKKoq2Rxfag7zNfWH+Sm0a/
2bLzGs6XTGuzNhdWh4T8/XZrTlQhpcv8yijqi6a5XQr1NbziQSLPczKK7IQ7PnjZ
zJat5czlpvRWBNS0mbdEu8KSPMlbaGI2fKaS6LcHGkFz1AY+g4c6qBJiR7xFYYer
PWeFZbcSbixS9/Rl5/vBUlTvZ9v8xyu0c0hwBExehyLTqs3T1tvYSFP4pYZeIv5g
2DH3cs/vDDyhecptQrpucRylatrPAutOEm9YYmCzQ9o13EPUpNwhJ5wYZHpT5wOV
x+0SPuuuf1bkrmfqjqta1HTHy+kOPm22ADRqKmJYlehl9RI6axnuQTVGistfOOPQ
xawFUwkhOjnDOJ7axmjKiHygUanIS6Yl9zHoiCbH464QZQ6kTkmQcHi9W1q+jlVS
c5eXKjuIwNKfGGHFXYQ6iu3UbxjcTlWG82nviDkeKiRFqms3Ybs1JZAUoLXSwMSM
Hm1QnRCO2EaE4FTQo0iHgYDsWs9GNKea9ANwL+Se93Xtw+u23LFSd/Zx/hTvkra8
uCJcexcXCf1ivklVzH8O/ALUl41WJLChTxn4oWAzucl2ETfHit/LSdlRCpXWliLb
QWMiJD+kP4nNoEk1ZniyYa381tmI451tiRL/R3YEn5yLfjICeT8ntF4OMzhnjnqM
iQR2h6JcUzZTRB//R29cTeGPmhgt/rvlAHI4Wsfiu/MOogEifws0ojgdlj3QJPbB
s8qaAD+1f1S974kQ+zPkxNcZW1tGQVEh73gzrWTdr83rO1ExxDmo3Zwl2Dfbouik
duxfvmhAzO53WiV2NACt0wXN/QVI51+GzG0rw0ikd6FVN1enUMV9bm43Pjz50zQC
FgU/2TKIRoMqEf0oSsgS/W9l/KNuTAEcA+9iCLKPaUFOMVkDtTng2ThOkykDDB+/
TkUqXEWAXuxO4rRpmlvQvhi+xSnxGm12GSBpgnQqhcDhCGXzppTZ5MtHgWsSrXma
s4pawEvvYlqaes1ZV5fs0w0MVkA0i5/iQF0L2h9H2oUkA3ohH9UnmV5K5hhoduyb
SmaWNAE5G7T6nay7Z5RmwL+ipJIwzE1ZAvs7y1oo7+Uq2Gf5VN0L/HybYVyF8gPc
WMIQVDuVjOVpWLxtkGD5hHNDrbJvxD48iQ3ZnDIE0ucNPAucGWzmS8u0YQEyX2AI
0W9S4x9kJhgI3a3A9gm3z4KplHukZ1c+xVw5Z3PdmCvaI4m39wSaTAV45hmD9Juk
3yi7DF3WOS3X2o360OdeHGmyzY7fwTwKt+TAS0lXikqhMb8nd955glSMO2Y4OZZ1
Tsr9XtxisGwkcUxzwx5E/VmQ1iKd8gHA1o3FGQiqvVISjoLqgtLNg1pD5VpoHf2s
lU4KUtWSk2zA5J8or08y6XdYXDKS3a75puvn5z+aaBcL3BHO3dONivs+wuCSWWTw
jsemfxmKmhrVWr9fyVyQOTaXL4GwMuELOE1HO1aHxi3HBlFkcJ8Ni8XvhRyMPYiq
iYK4VQRNy5oUlwQ/r1TjzB0z+LiAxS1usdVP+vHsTkYtnvLQ+tZQKXpIbQ+P0hEG
B45aQJl12u4zIcnN/8Jh4G9CXPSUNQPumXWufbbbW7q2XtmbvBmSOhwe4qYhuiP6
pticQc6Af+7zYIqWRPrKJJyijK+1h3GeL3Uid0P9LEemES65cX4HYdSQ2K4fHr52
GzalMkF/iIwKgz8rH3OyZOyK/OlByoG244vn3HDlZQjbiOPMOZ/UO6XCWDtlHzLm
yXdXHuIcPqxYk0E65z6MgIUs/xTiQON+JNA8glwm5vYulByJcn7+gKB0qq7F3KIh
Oo0tnHIcXGZmwZMZXBkdBBNUyx50bDet9TTrldEtFETfGj+EHVB1Mh79AFHASJF7
+EVlnUk8kA3+W87ZR0euta+B7eZz63DuE8HxpWZ53ncRMPC3gsYj8/q4Kw+0x5Gq
`pragma protect end_protected

`endif // `ifndef _VSL_SB_SV_


