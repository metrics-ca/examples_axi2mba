//----------------------------------------------------------------------
/**
 * @file vf_axi_mon.sv
 * @brief Defines VF AXI monitor interface handler class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_MON_HNDLR_SV_
`define _VF_AXI_MON_HNDLR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
lF7/192u6N7nTAweFaWgpflW54JhEbzQ5Btgoglo97N7H3d/kpIuEtmzwuFLXzKW
XibrrzavvLAwfdGLLONCQ9jHQ+Dab3Jez2s/IVBHL+gyXjli/iqqVLz4TqkYIRFz
Vwpip8n4/bVDG/eUPXXmOynO/I4DnmHCh+C8jH715iN45ZDXIVRx1/groiFH+eqk
c+Bo0TkNxh5DoJ3OCm51V2qdHBswlN9aehnSOPOMpPBjSRgU1qrexoZ2MCvKSgUf
C4fgjlDdtEjfJUEPiKSGRh2PKfzcJy79hVZihKx3EGnipockuKLOeoqPlzfGHJRy
6S+kUfqPsch5iw1/8phkMw==
`pragma protect data_block
AEakI9okLiH6te8sleBTMJLnXjR8EJ1S0wJYymbkxhQsOQM3r5rOzot2d6IecJep
Z88laCBwk3Jfum9quXDww4fB/dcnXTPpxHJ4D5FVZvb0aMf52q2iT9SV6pGA23eo
782+lWbvHXSm2fI83rDhwFd8Gr6Dv4Imt0FYnmLqg3AnBrmpd81Za7R0Fu1jtV/1
GILvExPcrBAdPejiGMwRpNk/HNju2hNn6TchGgT2C/QxwkaZuNgM+F4oqTTVDPQV
27oIZRq3IzLtc+l5S21+Bys53YzPzLbn75F81L6H9Vi3ndwNPfKHwoJ/uX68AJiW
HhWKs9LjeVwWYNvJqAsEknshzMyqZsAuO5hxT3d2dxkWnO9hbgFlgnP2bVlthM3L
eeGRCv+oqskCPgptx80P5/Occ1957E78es3wnShtQAK4g7tFDOAdsuFhRZUT8rAw
WriH45Kfo76FRffGMb5P7rIWY7qb9q7TFxdRwzhVoDOzLhmb46f+qynvk7SMfhKK
c6Xiyqj52Cha7RKDE8wTFgFUU1HS5d8mHneHNHSD23ffEb/DOk0xK6A/JdKFTXCD
zbNQFWypxVkx5j5vCpReWyCNyjy+yJbW23MgNKmwj3OoYkIur2nJnviQKdbCoUwX
C5c9GUn+dvA9q9YDZeVx5hacLClk1ri3oOq8PVU81R8Tx+ChFZPIuc+Va1fKTrAk
9o32M/J3kD0IXqRT4R1x6r1+UxMrD/sjxLAtz6P70RZ0UhEM0hJw/hqtMNdGFT2P
yf4QohR4dNS0KCABiJtKchX7k5deSlBfmh5lK3IcFpC6Ff1WXbDkO9HVGTOmnVk2
C310mU4U1gGsrqYQcP2B9maMJLj7HpJqxq90NjRHlrLQ2nWZMT5pquD+r036FeYl
jNQ6ud31r3lCHJVEBnTctEXlVbS869wjm5vUxmDHDtGzN1kLQt7C2octCUVlotKf
ys2XJurG6Eb6tlXxuiNfUekyZCiYuwjbAN4iLXtxurYdf3jDCQWF3wYOLlY3AoBT
gvlHcZiXQALcPozrVjBsA3Cc+m3jApwcXhyJbIES+9aKiplsiE92RBkkA+rZl1Xb
i3Qgr1bayizs/fa5JeDk0Gtip+WAaP9WALoPrnkEkxGp5q2zYknfcJTx+6M0UK+l
3+vjiW46Syoxsa7aqFToaxcoWS1No0xAChriPcCY57Uk0NquKmT/VMRRyhiFm/cj
uSFvt/Y4FEVZkL+HfgRT6zvL/1s3+PCgjcGLZ0HzJVf+1qm1YeXfWKXtTwsE0sud
NqSEzTg02Gpi1az2oTAAcIzdc1Jj6u164ogOY7JzWKdeQuKMPM6KGoQDMzM5P+G6
fPJsWjv33b/JVm339OUqHzRj5a0bFo2rxmNylfooqFscMRYQJxi8hsS3fa0SucK4
UBAHnYjveETK9a7S3LoKWIUuQolrywmGva5ybGwLv9Xr7KYF7PiNj2XIm8FUPTHg
lGic1prK+1exsqIGOwUc6jp2DhdbwmIUa5I+o6gAdBlKCu6Tco1jTMxK6Z+LQtSu
Gf8LGHKjE6uypp0ddbyGjzdyLCptrLhv0FTqmYed96pyydUxj4yD58fnCcB9wFIY
mG6cqSJzpFCPERy/r/5II8iGYeF182yl5CuHEYswL/WzDzQmfWDJqQpP2MqjGvSt
VHU72QNGf7TTgkx//EKFQF6F1cXOorcXp9SeDEGhUsgV+Occz+O0e7YLEE/16fMx
fg7/jXQk/wdF/d6KwkavWrFA2uN/NI6lDUzdaqxiRwnkn7l9kBaQxZX6TZcwafaW
Ur/NHrzzhId//5JfvjcKOcqagvlSRlXupNBPyUlnHd8DCfo35XoqonTpxHDW3QGs
/h5PZ1sYUe2LV9UMJmYyRgo32Z5Bmg4C0HjlusUs5kANnRa6icktjSTbml25UZTG
CCbmQH9hDhyJydftIKU5eDTqltqHPAuZq3cGQC2XpeD4Y8gOKDKXcGndZyY4JhI2
3tCLXj7s3WnYWTNnT4VrG/1Z+epwdxJ/2mIKATX4m4RPvJrLRcj2t30ckyBuIG91
4nqAbdcETIII8AWQxc9CJm2prxX4YWoXEjqGj2XRlvZxIyo4ZYWmy87iYRcGEfRj
uRz0hnn9wXxjCAPVJ3T63rh5QiAOwEoBMK/JOFrA+l2vEL1++5Y+StGAhyazffrg
wN8lzBDUZXVz7jGFHoD1PkbKMzeudIxDQDgI8jqYpsFJ3PP4N4dhFw0eBUqmKvMZ
wR96BX8df7KtB2lD/kEatSL3o2bTeFjgXGGObueYahancfB67j0G5B31q6OR4Hwf
gJHCmXQ98AhPoVtcoKxi4/oS0GVS+5cWYTSsMzP8fV3WuqJCnmnN7OEc0FPJDz0w
XNeR6Naspadz+mA2YbGgd2GRGgDUANY2SszzQUU/NjvqluPHoYm65gHVyVG/Tf4m
F3dm5OisSPVGb0lFDqDafCY0v7yjTk+87bAfO97MQeZ56iC1AVRr4fQze9MxQRAs
Xt5xbyC57DNxgH0SUb1vMr3Tvvw3Mdw9zBKf0wpG5mxM6etURAwRrEPnjHePK5Ia
gagKDcDTN5bX8Tc9RgmylD4Nb2PoIOkLpWqUxWRBzmdECV1lnI0Bewz4yq4870g7
gybn0u87/a3zeWXGebOEDT77yIBSDHYmkYZl6vQoX6HkUKv+iNALEpGxWNN+H/nV
X6kXe4TI01kS0CuKmqMpo/GP4jTnh6bOihtm9scc5j2Zv7oXzpqc5uhEAkWDcSJ3
M3kUXK1Odwyy0cVn5hwR75nFR0Te4SrNFgi3ETR70JMQbi81J6XAOhuSyVT32NE9
1vnEYXgin/hO6kHEXC6u1a+URt5z6PwHaF9xdxUDq9/BVswMQQt3+siEy3ElWeDi
HXS9ja26OslM4yKB+To3XmCbsSo54fsKT2cHgj3AKj0p+9kOOekFo0FsBe2K2YAq
suAQ/ivgf3RaVL9ymLCIjzfeTKe5dRTM234vdJXp1+q9KpPuy2vkV3MMpP0sAX/I
4Z+iABXJ82vnl9qNYzmBexCovrM/tiVPFu+6V7/mAswlCK0zmYO0SNF11kjlLXC7
BVMzt1h+8FXy9Uopr+3/w0IVVMjzukyIIQlmPiZDVGMkwf6JvPhnbD8URsDoOSin
AIirWB86ajac8QG0jOx3tLlL94qwcYipJ8x38fBk4pzmJxbtda/Gij7HJMdqydT4
/2Ag82mMqLRobom32bTTPKtH01s1VkwjyF1wDoLt8LFeGHcSFWSeKKkR1mljAzDq
Gs+PJriYJoNUcMytomCynr2j1xpDqtMN3sF2BszuH1xRVU5N/7NAfFAq2pXF5Npr
5tiq69uHCFQWXspdJSkiYbaFrgm2vNZWu2Ia24OYZRhxlbti5OlLfx4m3frNSl+U
yzd2Mg2o2ti3K0PSyIf+DSFQGM0wA1w2jPyrFdynn+gxBM5TexCYPApRp9sHjhoC
KJbFPGyxVSZh1fqKoQc9HrnqxMjD5mX06/Qb7GXyT/q6swdlzZa9e+c+6Z4xAYDt
5hSN/LfMeofN6sk02gdFptK7wJSAuPuObHBQyHjItptH3AXr1xpNrwyNNSZmyL+e
5PYY4uyrX9f+fLwAaBkGKdVCMUHBoS0t0CvOAgHWhWWvWcQW+3YkuZCRrGYjUAQ2
DVExhdiHj9a1Ebwgg6Aa7kyQoUJyKF/7j7T0vAsGV0MGt8CBhcaURQ1LE0DdXDph
kZGSnfUi6x2Bicd4MfswvwSXS7gJDCCL2j2+rSd1keux6h7zX5nZ+yKHHDXkS7dB
DbiHrqw6p8UahJcZ4XM0Tj/C0vBlVZWtdF2dy/wXPwpNFX3MHdv5Qzug4kjGfBbi
f2iwWx+lTIkfUEPREjjX1cgV8PJhydZFOxXi0EeglXTy5aLG/y1flfvhgKbuuqnr
f0riUWOyjbS9VUA/nAvBHqmWsHh6XpWT613kJyynmBDRrpJ2oph8FmjsKUeufg+f
UGTj/6poYRysrfuFro0y/wjSEIM66T5zGMXGZpanRnuxT7JfArSWQx1XPDUCa+Cz
IumfY5Wj3pm7Ic2jlHmuWzX5TzA9QQ6OgiTNraoyYF7vVGZUAd3xBw2ymUPlmf8O
mZXKrOvBNSSuS+WmV+31qu2ra7pYmW0qZH6i9Lo/muCzs5dyV0CNJOlZY6UcRck2
YV08XBaH3P6bzYb7TkqkcTkL5uauKyGeEye4I4/JK2tSNFrqZZuMUlwFAhdGpSQc
b6jzeCTWTbkAaJ3v0Pq88p+bAVxIRu3W7XHpk5aUXCtQZlyNoUkehWJAHe/DbjsF
6EAQ/n+hmpoyp+RJYdKWX3SN3GfAkponndnQ5QnCahtgrab741h/CEFsdCqYXNnQ
dSJDhRvKJABEWkryh7J1tYZAw0q8r7DmtJN71itu3Ywi6H3fySrQv7HX6aPCz7vG
jowhVyMm82JtpUun5xuC/GoR4k3jSNQevNmrnOAOcXozjyKBu27BscwLXrCv8yPm
J8ESLjOzA2Uc1/FboJAcW6VH2EoiQJg026ukNeQAJENfxvtYz2lDaP138AjAm4C3
fPLPntshzRhNAdyCc29fTztT/YPtn5+ys7y9f04ddRPHpJwYb4i2/lqkVkyqIa0e
dbzFJ7327edZszgrpn8AqPKBwkZd3Le3LD63VnIYnqiI3aNqEiG5U1NjMSIgzUHu
+pBAlsXKl7ZIWpOk80aZ/+MxRVGknM+WcCFqe1RT1J92xsmeMX9qAEZmqDZehAyc
+0xAKIcvURql7TkZqJUWVEQjOv9kmFayzqUFxNfGcG+XKZnwr97WGBS/4cCNq4Pn
QEJLkaqtgmCQN+88h271Pi6VPwVsKtyhTMt/lJka0LfivI9jmF4WqCJSVM+G5qtA
EKTuYYD5HiRXf49PHyVx7majUnz8BNqbIQahpN0ufHnBXpnHPFD4RKtdzZ0xfyl8
Vo5km15c1Phg71S3Zea/mbDkg3kXlpile6Z5XbM72f+KHEzSK33oz2cjT6KrcmyI
Reaf5G9CmelM+WbMEKBIjm/H0ORtl7eGICuM+INDhwOycp8BB+1SQQ3iquttilUV
LO5H5GJMtf7AcaVzu1hrpSP2VhI9Z6yfScPLBqS07a/DeeNZu2YnDeMoa2CTcY14
vyYMEN4vZhxYT0mZVBDl8sjc/qQXYLqtM2pwBL8fut0ovHF3gIi9axWAMbZyriTy
pWq9rDnIHZBjqtcE7qlL3bVDofq8sWW+us87CjrpouIJWNiANRgR3AzwPxVIiCPU
83Mvo33qAQcgC12FWIwBL0RRWFoMUFjsE/7qjVrlJzKddrQ+Qe5Z2Nyy/g4Xly7O
H/MQhdRJo6cCh++E1LnYAeHJQ/+nUJJKYjTWOoWicbHoHzl1Yty5LxwAzMkQKGB8
DRj7u8y0zZNRL2EIGYlhztmrU7iAVmenS7aDaSrBeV9MpHWeyc7Y9tF+zUWMaoUJ
kmR6dQrcKMJfF9m5QKv2ngMOSX2PR8Ft0RLqPd5hQwArghIO0y+qcAatKY2Jti7k
YSMbUorZ4tDHRIuXPTRsR6H3wJ9FPzHZB4W52gwlvabsOygDY1AemSiifDtB9etG
20plN4/ceL9b4smiA7zRCv38dfA814BSDva/oYWd88Ns0GumcxGZedXITE9iNopb
7W1ns3t5dav+WpkqeYIFDjcSZVNmJCwo1ViCsx/bD6M+9NFww8RINDOd4YXdgXfR
B1VYwVOvVZjUD146tWNkGoHj5tnWcPuUTipA/CEK9mGfMIPnLFxnjGMT6k7itGFU
WDb63PV4UGqKreVz8jLf7H1YHk9Kvm9ermPmkwhcDSWLaeNZLVfblGR7ki1IRE0L
is2gAdke0E5BmyD2NfhgZO8yv1eOrTLbLTh8fha5Pmzjx9IoPDx3MBiUSRnUhHWs
GrBKa0kRpJV7d6VSExQpHADm2uTJW+kx0C3IkPkwKFxV2M3RpBsfttQPUT9LGd7i
lD0YnJ1rAx4uxY3+kzriCjTlX90m1J9w5sMI+wStx1P98SB/j6wl73oF8AHmYiYm
EgPSNQGOzgdaa8oyfPAF8nTw4xM/IBICa5xqFzyjaiUvTpI7tQOotkGs1S2KEuLI
hw2Ihl6+ts++zIxLnXejD51kGs+JeN3n/H2l8p1NSivep87gAgyCb5woStgzr7cg
ROQtyjtuBFt8haah97lgWdzcWgkOs80bzGXLXbixgwmDw5g98DZr7FJc47osqcmX
aikLddAIMNL0ZBCHCRnAg7yU/5K5UahAyzqOev8zjWf4P9Xqqv9fI0ROzIQxKQPO
3bBSo9O0enCLLrZZeGxzrSk+LhWAiQUOmyhz4STZjDfYYmO/RYPcJESykxEZkhjz
RKHuWq4Gglzs/ukll2CzjeYY+t4oYhDj6FVolQRO5I46IrT5qDkMCqu9b9IIBm+B
a22Mp2xhg7r5llv0eIE7SoRznPQxFa4qyn9gKbH7Cacioc4dVRZqtfpwjr0AeSA3
eAneOjp9YN537M/3D4EwqQkeNOtPDCsyEo0bQieuy2A4mVEYrsFnw+aOrg+NyNcR
5WKXz/kcP9Te6XKm3nGrVK/9XdJG8XDk2Vl60olmPyMWgJJVccXIdTIIgVHg6Kny
nUr64lT3sIvysFnw1JV82+S4vf6HNXFkMaxzIcW7tJEP6Va3fFjf+i8D+Huc5SIz
fr0CjLMzj29EldvnxdpwIxqfTTi2qRqyk0l+JzTVBlfktsuWWLs7ZKXUwbpqiX0a
uoFsXspEhrGoRXLDCzDMFd7tNjutjocr311GbVeacOfr+4Apsl+FAxrvrk+W9bQy
plhJL1WJ37kGHSvEzaDwqaTR1QhrWpJ4vmXwKVkWkLRCkRPjVfIDf1U74isboi/Y
trCLV7Jy7U1nGyj8TCPhX/8A5GFzIImQKqb4H0nJQkZvfhlifXKTxChcBSkM0wJd
el7vx6f+dn0daJxONJtoF5UFf+mboQSA96AdSCiGtFqruAIgRcNq54aIj8xBur1Q
WseDnFV0g+OLE9EpeIvNxnfK8ERTq7cBMdGHQNOy8N1clmthi/OVwF3HfLAfhmGU
hksbnRrmHXfdKKKquFqkijg/6THNRMl9TaMthsNL2wP4dhw41etfNjOvMF4RFVsJ
2zKSmx9A4RfBG2iusa5wNCzkPjXxFICj4WqJ0T00U6TR1wDtkWLNWfreaxFyX7Z9
V7OQNaM/KAQfUir6B4mbIIQtGuDeQ/kthpHSgQdAD4P9RWFP3kMhFj5ikxonsvZe
L2UnQLa+7XGbw0ybKBwpW7JLWzdJc2JWL4zEJDhl32EsYZ54sAgR4dlKaJlU0m9d
4KjrH58mjfbhJwzXv7qYVJQvLkYQw0SrnDe33I2Q7HqJSBdJO7ioGewModeeNnD+
JaLEnybbu0T+z/WClHeeC1jfx94rur1RVAygnuJkEaUUF/RFIZMlIvsIJJJWyXdW
j0judporqd8mTRLSHdRuk+EiqLOuS684S9c4jT+nol5HdoWn8TndmDsXcxDqjr16
IpK0cQDDXx8zUOSl6Awf4IMRJwgwONhyghgz1qETAJKHBOgsCa6Rnclsl8Thinky
Z0bIQRHpxfjBQsvmUkhko/5AiQujuQu0ryn/S+MGRduUUXrlaKY5qpw8YF5BF4Vw
G2A068XOciNz9sXZA83/So1oJZPuUFYmATO/bT3YpyFwZl3q7BlGHXG7N24hcsHY
UsIDiAok7xDs35hCZw2pvP6ATYSzdqNfbe87bqY9yOdlJcKU5WXLNmT5xra3ABjt
k8pY+f3rIInUeydSESXkDrPm3jvNwKStm6dyzFh9bhP444INITpQ1aDqf1ydihGx
WkerVbuba/5m4cE68RsO+/4Y0udh06/CM9yryT0JDvmOdMkK03WpmfRgSHt1C3tQ
Fv5h2zH/6vTKnQ+stt1or/9cE1NQQrYeFtoXp3eScCsGYbaayIjxZRYxo/IcDMHk
rdUoulAr7QZzrP9+3YHR4rpjNEcZMLsQBTFL0YzEETS8M6BnO+/+FoglQORKDWlx
7gw6HruTG9RtzdLXFam28pmKkHjyFHPBNBjTKNI9BuI3dFs7y4M13n4p3z6fY5Hg
I/EKmMZ+S6THuRjtohmgl2/s7/2Gcx56C2zfEfz0ltQfdPwYf9QiZvhpVSAdx3RY
S6yQ0urSn4aDn5IPX6ljTfhCyqrk4PYwYU3DOZcJUkpBU0EneB9ctNRX0FMAUj6A
NbCAYoz5jheDUDZ5VPSsqMDum6W9rRcYalPbl0dUYdIsC04rh5ggG7/15kljMtKI
YsWLNpEhMPnHIUF7PmOrB8fpAbgwivf8ryXc5yQeW5GLfR/fHJ7q6kLHaCqZ8fDG
vmo8rKR1xd3zOppWnlvqFcxEeH4lAUVTxNh+UORXxsv8tpdFKYpYVP1igDdaU9LP
nWqMi+eje+7JYRTh1YA0wbTS3MXdlyqJEfCm9gRSBhn0YXxcsl3w649LNgMS+F1W
qUV5aWk6fSanR/227BkXK6/XKabLNUh6SYi+N4wJwOkX4dMtcnPPtREN7uZUaAGW
F1PkV4SV8BVTDrpuzuW88YHKovEGbQvB8FmnoiacRwHSiWxkuSaiVvO3qI2gHK6a
2o4HZTwC7OI/qz/CFnnBMx2czZILWrys9//EoLHtDJqtXOpIFTcxTV8MkHRO16Bi
lALs0QoMn/JTYdUiSYJ0Rg4vA8EnunF3s09AMVgJm/+WGJugbBtgz0ke+jQ8+Cy6
MnsfWyXymVcDBIZgfW8fb3Pe6glzYL4yVkfFyE6hrUz+1awxZMh1EVCvV6IuC+4m
vtZ4zH2JJt3WA5XVeymmW6dRR4jvZVHS3AxVTW/+abQSwI4rJWqWP7rQgdI76MLy
dtez7jTXlY8GpiDjhtkb2jHqSVPbXBl3sFuQnGPquMrvbqGhQrl1kflOYxBCsMrq
TPCa6hdY2PgaF3PVUPVV9sSFFY1Sg2+qhuTUWgI/a4aPHbzu4VsaIzeVZpAwJIt4
yk1eWBoqt6O2D5tWz46GtShzkl5VjrO+ne0v6qz8gbcWRYiXcv4HU/TtbCF4gc08
/p0U6Hjj+Xw/+oxMqkipnuCZDpAbQN56NoCLNc1EJD1Y6Vmmh79+g3VBmFUhAU1W
w6Cg7hKe3Lcs6AFElQ5Rttqb1Qa2PvU+jw6a8NKddbpf7R3dcUbCjAs5R6R+3g0e
DsLmI9UY5Kf/nmGsnuymZCSHCTmTOBEAF//LLTFOSqlWGjpwkRoQidSLI9Dl95Jm
MCIyfeGo81MHxmQXd7XRU7WQ76tps1szVf9WSVX4wuOGbkKriiiZC+i2hGAZf4Qa
8jK9sKO/oGRmLwY72g1AWp4hjMLD5iOjzMnXnmCHTWPD1rARlKPxT+vBWqCsWnXI
QeJJ106F/Bkfx9nzG0Q6YkeSkymoqqj2QA10eXGFQD5BuLseFyW3qvw5oUJQiMTc
OKq5Sk8dv07L1ft/Zm6Q7P9Jskh+OksC3QCye4l03vDTsV3XNlYucE6YmzdXYjrm
xS70WGEkh/hmEnXCj6Ij8zgJx18q3N3nddiWHjIO/y4kDexv6oLwJ7xdVckj6g4X
iFkjcTQuxvb14xr/pBHHAv66ln09ZmmjFBczHivadN7Fts/bFRY5tlTvnVu6xNZp
0qLoctnzOSAvTi/3eESaqQg0kQCGo8UxU2XSe6J23u2H1+wEl88hd2IUlAaXT44G
XHm2B5yQ8jBZcNI3WZr0WkgrUq55kcJ0lUv2Dusz5320ICeWX/Fum8eo1NyxG0jX
1KyvQSMbxOwq1FbzBI7FE6fWzVM7kWnpJMFMbBNFRziIdaA4gAiLq4PZztx4Iz3g
a+wLQJ2CxY0fzjewWr2eF9mBC+o66SBsMGcY0JYpD654VQD7KJ1NT5kbCXhSXQh0
CmxxqfFGMpRzyBC4Yg6eTL4qwkerUkEmvMkhEp4++Fb/egU9hXvFHi4o7b7jFWxj
OuiZ9xiiPQXRyCJuP8inRHnlw7gNw7IWOe5v24XWtZy/ZU1CTTF26WPf602j2kUB
G7y6SXFnVtYIXLbLartf7Q1LvRvFWNYL7RWlPsxkqrDPGGhVe+Fc/Taor1tm2+WM
VqusauVhWbNdrkP2phHpOs6iuqNW4atxCLt5wCO3snnMba+SCAjj4Bv4BmS03yJD
gz+bTHjWObVvSPfY8GCzZsG92CXOxjAjz4brkDk70pVRumoL6zLdY3MC0u4DYnAS
qVQyuTcQaeVcbGXBAc5qTI1f8uCdigHHjRDkjj3tJyGa3kwdG7PKyiZnvyiLxMmY
SCPrOerZ9XdABHBkgQ+O0P+/CO95Q+NA0eqfrtNmZafne0Vl2u9RvvY56+xlO2mJ
T5acq2R2ZjJfkwUapLvnISzH0VD8ON8DiMbwz+EeyVFDiy895k72A2Bgpzhy+k0u
JWjB7CqiE/yzlhoVmbOFLJKDBWySk8/O5xAQXRG59yPa9hARNBgyE6iLqhTEmuy0
X72CL2GajMxohWuBWd4hcMr197NvBBmEF+YN9c9KnXGQsGkueE08DTNT4QR4HhjH
F3E9DEBpfaFdQWa0Nc2fJ2JiGyhZLKHD6r/N3ZPzL7t5HN3kDeC9Y11KRAGT9X7K
jyH/DcMcZV9+eTVSsuHxSnCeODWskl/uCj7oh9/P9erZRbqpE6O0tQBsz61OV9mI
8qUj+aBe/MaaX0h6C63VjXZThvS3aOCbv6Lstrtb4cVHjuvEt1tk9aceShnQsI1l
QbBmbp1FR/ByjN6bURW+oRnDX2msSx9YFYD5K38I+x9USaCJi0iGsKFQBr2PBfhh
SFBO5wzlMhaRnMT3X2Fsqvn4NIvE8w14fvTGtPX+uH6qXFVHYEJMYgP1jQ/m0kIi
lT01uSTOwmgxSIyKbJHpwQHi2UK3Oce8cBR99H0arZYoDBaiLn8rxjMt6+5goVie
SxITabVYvpuRp2d/Fq//XHQwVmUcDd8p6pMb1VbPoo3QrpMHn/LqGpQr1p119nnm
3L0RDFrwhaqdGRJQjBLtmAeDQQ0YIZV1KCoJWd1Lh/hiHtwWkI1AynXV1oxviiuJ
vkyJ7gGHbWCJKO13LbVQ8JnkMQLPdjc8vfMvVtfSaS0CNZYWq2PmWWMlp33LEheQ
H2sOYo3rj8rpJQ8QfDv+pkrVBaEhyC+KZe12cWFoe66kzb8A8PyBbCzknmSGcaRs
dFhdlOaA3mk18zviB23hB5Y7vEYo2y+9DoSDAwqWIHc5hq0rrIlBAaRGZfCPtqnj
aRvfB49PCOzFKJqL7Yx/E/jeVYRzvRq0u9ORpAQQSQYCnY8H30GuXT5DuUQmNQ2V
CJbsL94iXiIFbPMKfPJNGQV9ux4tfSxMM/7eg/INl1vqH2K2zeAUHGJAY8rhI/Dt
h92uNFgNYhvEGi+IAQUE16Bu3xKUk16yiCbv3a1yA/OG3BurH1Z+T8ny6EMBSsrN
SVVo8rNNNJoKk2WqRKukrhZO7gcEUKJ34/lKhu3DORgZm6o8jSUX3XIQPoW6TxqF
55Nh6l0Rzd14gD0vX1pFA6P61P/IBrxFiRedw+oBy9fCBvmLozTz61UJIqVCYpma
7QGJE7fmnJcEc4SPRdKys7wxdM+ZdlxOTQRV4p1HpazY0sNJBU7t68fOqrJAh+hf
jVMBZN/y0tSedK68tuNylEof5KKojE8RSLd8pxmZ8Td/s2ZSZOJnfL7/3gT6SysM
aSDYadfHMlToglzJbNSVvW56yuQiaeHKTsPhPGJro/hqmtRz1pyYG21noYDmk93g
IPl2UtIcSM9p248ic/GYn4ANpKrbyPbQLVpZguw7NlR/LhyIe18Efb6Asdq5ji5U
TgH5NDT/EVznv2i3wQGTumYo06XunwgRzP6OS7LRFMgosotcBPQottprpRnChUSF
Pr6r9x3n2DpQUJ7subkkhTCSWXjOIx7JKyFqNSDU3eCgqnbelF1SwMtYd2jj65Us
WL83nl+y3IT7cIZmpI/tBrafygEKbrRyctZHQFf1vNYaUAg2j5q61PpPuc2JKJU5
nj2sMp52r/d7qONBI31DFcXt6uy2GAKcFgA5paeZf3120VhyWzz5VNvj9FJgcB3Q
d2552XXjB0zvvmjOHfhGD/1AVCijAwbcd9qnaUKagmdqgrn+EKE2VXO7YYdVK18z
txXkpGYPnAb1r1JSsiRaSKK+nTCMiysmRhI5gG1GdCEwN2owPw1n7lPgveIllyP2
r0XHZUgnffEY1K45hzotze7pdzK7pHFcxVlaxAPkMdxKMGvUld7f25txcH9HSdvG
KKZbDlix8PmN23m1mZf8EK4AZZw4nggv8F8I04tNMvMeqlWn8QCXjnQ4LEzNE5cT
DUAbDQdqpkpjnbOH8gbZ2n7W3h1U8PQV/Hww2g19GCx7X0woM/CIFavNbX5AdNVh
RdLgv6BrLBl+iNyMiolH7xBIkjpzSqAbvJHyqLzXXnVc2ESmDojOeYrIuTatOhfl
X09H0tQhxUXcyDWCvgtr8sug4lsyYa48+Eu6xMReKFraHY3tnm8eB1iLiMxrjNQg
YbJijt16Pslm/pcPHhnmKZoERdN6cdYLaQmLi/1rscDrT/ATx0FmuZ0BFpud3T/x
PtYSzQLIZbTXFhd4Uq6z883qCK87sHVIQCJgEwwH1uG9oszzXgtG8ES6/ks5blO+
GRL1mIQ67a0PEUwQjScrvGhnr2miTbvrrxFeEfsA7goO8FTngvTiJ6KWqOiRFQm2
v2l21aznqPIQRt9gKKdhJEJoATSUleA04r+Fpm68TZrSdSz8jt2MRyvtD2W2YdIF
RzVw1O/ZL3k5aw+BMG7Rn0vLBM494V94hIjtriRQ27YBapGwHOMraBSTzZ4TVUmA
T0omluwwJqZByWyqNQrrE2pHubNBNMIJ0BbcI+BgPs2/2Zo99TuMj2XaIaSxURE5
ScozkiBodjCFpvcDXNy12uBPncGBVKF3rAcbZraePwCqovCwRdaZ5411h6IKAKfE
yPPITtCtLh2K7UtNNSvG8YpQd9zN+NGK8iHLxWWe0KIKkJQ1jp3NpXRC7hR4lmPy
YJwle8k/D/8oDvqeqaVG5Il5ECCQWOBJkVvMZcuxmXnyWfhBk/X0OhVnt0OVfMk9
7hRLFA4Vw6K/twcjWKVShlcOvGcZvT0ErRIrXzLrPs4yMZEBPAlMOaXpDiHYsd4i
9IkYxNx7zj+wYhgyjA1AA04wdItWIC34g25lUrQb8KtGovGEcsTHT9k4Frwb7nck
zsjcqF2HX6LD3GaO/T4S4Fw1OqUC8OuM8LrBkIBDo82iDm0wLDWXg7hHWSuKRMHQ
iBcagyuBUtEtQPFER94+73nM1dQ0B1p8eKUD48imgJivMgxd/59zAvh9/RtyK24w
c7wxtQMBnemDjt8zbqeZFYWgj2aXYwRNiKE3ZT4FvvdvJax+VsP69OyPLHmfihmn
RqfkWHCiCoEqzUOXoDyifz0cYHeoev7lDa1BemX7iToIezgQFmCjN7DRrmN2vBac
PsaAeYF2D0lViuAiMitHKd51kj+r/LLjzlKIp0o4rNBiNLC8A1xCUIqGKiWqhjvB
X5HRrlzGPAi4g/dTpfYgy2b8d/WNHv/6dT3EJQqIXj1NDf025QtqPeJ9cvjEErka
pBydREJupFbZnmPR3PZMKLRNniwf05UTzTjC+GwjRbBzdYh16a8qnUY2O3hleCdn
/pPw3rKMFRoEE2sPG+wVVGaccjaqwGAmFuQP1rHaTMse1nn7wm8Jge55/yBPWqA+
+kaPpZtpKVnEg7rMInIAUCVUiuc5rLgbWYsRlIh6663zOiD594m+bUS7J5Ri4BOa
bOFVrpd85OP2V2P65rlocCd53XCSOJkp5XKeIQVnhQST73WWTe1n5rmJSg3CHXfN
o5WPv+DW9BpX7EiXKjtJX6Qciws7vD9aFdx/vu9rU3jIhK0nFvj6G27FFQv6tJ37
SLrT8vEC1ouEr8ckYIW9ckdz7HAemAgoa1Exkp2RG96HOnSxqgJISEZj4bYBkGaD
xLiBYSgH5NSG0f9icXgXIju+zaAC2vnveSwUYKnTpz520nIKtQgG5/ymokuSFmqF
nNg87svyqBH8p2NjmhswEn84dhUFsKLZV8pLuuA5i+2Vu1kqLH/hD1f06OvJmGw/
GV96d9j6B5rrnmeXzAUQpg9VEshDU4UA6S+YfDA14VkqNXCh54Uwqp92VYK7X45b
ZU+F1PybUqmHA4hMuX0vbz7rC60XeGoDoToNdnXBbKIgVbHEC7pC+PBphRQ9H/5F
ObLHQ6JzpZxPW659L6SypeAPSnjMrK1vm3jlZp7uEyu/1GhyPQSWAbYN51WIGi+C
6aaWDQlmFN9ChSuAl4qHgyU1SoSokXlkIWIWIiRjodRLZ+QNpxT4XhAXD7IQxK6M
2Xxbpe5tY7Alnd/g0tYiydXcKJI0jvWAZeKBmfVoAvZv/6o8EMxCfY8KmAQMLGK2
Z9fA17arNzmuKdWtY4Lw+iSotvFkjbwcirB3G+iBlMqLC+0L0JQ4DHReP4Tj3miZ
XLfgiN2KXrkWjXlvAujXBS3uo1g4v/SEWTafCO9n9ymQjLyGuZSi+WgoVleWFHN7
wWqIEHYNEll8r6IxCWwe5bKbVYkEOhDf9/cgM+mOAbdnxEKme7cRStXKKUlBbUpR
3Z8NQlZfR+M5kvWsSivDpZ/igrkkb4OSNAcnJbJ1OykStfVNfgNBniOFDFa+eiVT
el1VNtrqTHoPt1x53elKBTXcUbV6WwU48G+petqhBDbH5KSdOY2FvWzT+61ohYag
0NPJyV0bcLV8iMETLwIAQDvqSTzPeXWnp2bp/s9uXCfie+uRIo0EkIrImrlf+BO4
Dp4t4Am/PoSuD23p7b4RQTCeHCUjbriS5jJsykeLkufuGUp5C8AmUE/LbTyRpU6A
Vb+RcJWY/fb/I8CZJuTpJZYzWXH/T0aHcSnA2UTM7i9o7PE0wxZllM3DMn0KxHII
oc6Njtkr++UqUM3m+0YQenkzYZ0w/RWRCpq/PEbS1qAvJUWoB5LaRoRi6PVOBqXC
1SRfvLEKV+kg+JqeqZGbjAcrheOSq6997Iodf6seft8T326ilsEzbX1itcgUroVB
LtW7dDoByitvf5zKdi1KhRMPCFN3E9SNzo26UE1B/NNeIPEfR6x4j//aEDoxdwL5
TQsrdYCZoTxZqpu05Ow4bTCZOfW3H3+iRnV6y7VEsVBa1PZz1ceazRWPuL5xxilE
gfGoPuAgNy6rUcNkt1G4MKX9NyNS2xPW9oazUIQFh0HjA97iC+78P3FkK/Cq07k9
3YSGqE98hpEL2ZXwsEbOJBgdlGplrgi3unGqYrDmtDvjIkBy4d5ErurWHRMkt11G
B9inJVMhRbfD4qXBywvd+WUlOZ7SX6lYKYuvRwxU5AbAC2nKV10zuWk4NxuyPLhT
lV6MaoxYm15CljutjFI19oHCBYuUl8zHKRoV+DRw61JAKMw+8Q8IxPmxGxMXY37B
xQF8ewKQJjq0jz5rzBdW5PNy5Gt33WjRNRtt+Ff05jVascOgA+sX7ZrbBxUIljzy
JUxBy9VSsijggT7sE+T0rYK0FYFrr129t2WXjx0k/NOLnoGAJsi3ujgn3MYlY1bM
KPL43KdlPKfOlH7aLSEoyiYibAdRy04s8H4WAc5+EKHBjoxFmQfLFI9qyN43vbZD
vZxTSsceXyx2DTj5a/gNjP83wWsVsin4+5hfT9cyLKudjdlI6G9cpS6KUi8ScahB
IHS6sTAwkzIwjzYsKlsk8qyt5w/2QK43i8AcApm+tCu0m9pXMKd1cl8gfTA3kEAC
B3LHoAHgaWgaHe30P2xurbpmfbiLih/R6g1GgSeC0//RXh3pgvOmeZpdmERsHFwI
ki+0LE+iNb32t6e5Oa1hBtI9xd7swW6j9cul3dONrpMUb+vQ4Pg3seepCShaVA8H
u+WoHFUsJ9eHTj4e1OAlmEaMlQETyVBejZRVwf+xMjGWEYiKMZ6ygu9W4LQ2JaUF
XmBoQP47gjDhBcGtPDcmqjsz82IaVsgKEQEVgxEzuXRNhrNRnI/K7JfiSRgbDFZa
MOP2jpxyoPmvKljFWjY3uGNOU22TgVGq8rmeDhlA+NsLyUlf96DyMqaS8hIdsXOO
duqgy3YFChbG3klhUarwZnoDk6YoZCd+mHI9MiDsJcEyq08khpg3Qgi1mJRoiFOG
RXENNMKZ6lHa3hEcq5EEaUtCU1HuKaB236h/TUq3GQ3rrGlbniIbysSRmYzbKuii
iOH2DfnpH2fRhSrHBRppf+XesxxkHvIv3mdbuoxfe7zHPi4sqxwiHEYbk6feRdRZ
KDgqEkG08N65uMTQi9aXt+fLMg3fUNwzp/hAU2ZIjtnLzNYbkI6RzqcTANqs5xfE
m6+1SMyrVbmci2vs9WrpVgMrQ2OOtV8KDKEljzrZKivLR/k0J19KNNLzTdhIj53/
H6QrA9W/8/VgzR58uHFK8PfKZtsQzQHfNXtbx2qHFkmAobyBBbaBmWushmLTH0Ug
Z7hwcvQtiTXyQS8BTtTsnWVO+QR5ppekzRRenTlHBjRczto7M92z9/z1ekq5vXWt
kOhGrcafAFv3xWiVNB1hEZ/kuil4rT6A/202ZidVVKSHeVBcorsxHlUmkayNlS7X
1fpYkXsLhiUBj9d5hThOTIZaw5dPmQYuwxVBly5A+uRNRbI+UCmO8XWZKtvL+A34
D86XayFeuMBc5IOQfBUX0OJLFwB3SvWk1zu8VgZFjr1rBBCXlLpLyamU8O7ClOYf
nJj5Oxyj+HB1D9tLskLDLWKph6wLL/JC0lgVEabdlZLCgBdlgRc1AUiASn6R9FMb
cBBj+5FgC7RjWgRGpqRUfC3cbIyI4RSN5xceS+tfW1b4J+L3Od27BR6L65l589TX
OqZuZPfpJLqN/KIhh9xWwQ6blNaBhfx4If/58FAI0WbXequRNqsG/w2IoptCuIBK
/Ky4Lv70GFWeUopX9lY2picP7oSkENGlyrt5f5sInS1JIdkSbddepjtSePzt91n5
OxmFu9xyMiCjdIAoXZEJH81DwyvrEh5cpZdsb5mNPzJReT7rVuEQYYeKxjUUuPaw
H6tpwv4Q6+KQ0DXvnGbHRpmVZNb1cfhAVfREGyEuE3QX8vpSUSURZ3g+Hx3LGlvW
nXXpYQ24RwqaJ83ZJdo9T2iu38A+crzpzjTvi1c+iKlZ450VWF+r1g62eiZcm2fg
1njJwJ9+kw9gHMHmLaqDWPeSE+HYa2wKpdZege+AbVomY1WnKurAt6XocOFrF1UJ
UxdXFgRzsf1BiBsUjDDaexKQACIXuplxRez1m19NcFq+ZH+ZtebxmT2poW/YuzGJ
rdY44bUBGIKakzG8/gxvCmD5PCpUn+PDGRGmzQ0WVYi6iPidzSTJU9mS7dQv1ft5
vPrCiw9iAB/8Rlrpbe2l0wJihPHGKJcr/WSMoVeMWq5lWxtraHvRezXtLN0vST4q
2XjJzxxzrGYLS3Snx+TefO52mhXkBXPR+4POCCxPouOKhH3ZvpMpyvwEI2axTrZR
ktb8JzIqo5seiG+YM+7BnBYwNA4IG4appPQ1xMtQUdgn7tlMxFJ8vX8BZb+Q46SN
KQAeWrlFIzNuBbTGm2nvfuMzwmMSNIi7tykdAHcSAM/wYJf0c/Na7VCFHNUk5pdK
ViGpkKnxBhmLTITmU5YSfogTEmYe8xNrcq1HsdFb7xTI9CwIA5hvaHqM8/Gaej8o
b3llCJYBymmJjGV5PgMK1E+fjQG32AjpS62Mreqp+9HubDjtrUylHCZAyoxRUgWi
YFWjjBa2G5kUSKrz7ygAkveiYG+k8ly1n3nxuqZlIGhq7tTmJLlDwf4uoy1OZEMi
HkUiD1elGt1SHD6w5aki38DUBrr7eLxDSeS4kn41sc+p41a6ylzqP0t4RumTLnmN
j2tuLMy9LUHy8Vsq1fgk6RUBHTFFvCXgdkfKoYxFamHIn6yvyyW/eRTKLZviYNL7
HzrSwWS6TPWWEhRBHXDaFRHlbhVmoBbyiVcZwp9tE5VQR9zdp/JS26r/HT4Gk4CX
/v2NQhPHeFKzUlZsBuaIO6ZUrgLi3WwPe00+lmj+a4pix2jPobSjfnbpT41Bttvx
BNioQ7nOe5tjt0MZJ4t+sLDecn7xD5oXc534woP6rv/cGNOofpgFZBXBXylp/Q+V
4SUGVyGuT65tpp72HYegS1PnMJE8G3e/ZoOfXkPkhNqHIJs0YC94ylzFmsuw3Dzo
Lw25Qb08dez/BAKRIKlmp5gIAJU6sR4uhtziuZrafZ0Gi0Ijo6R8ZN9EyAx+7hXc
mBFpSDsdRBpBgA+zZl09F0xt2x7KDuY8f+VoI3OqIVSS0VDUsMly43/Uz1jApvGn
SnjQEvoj4cyXIRq1H5PmUUMZAxnfC40Te/k4h+tRpT54SP0FEF6PTFBA1HAy/ere
+wHkxaPOvpn9kcspCIUKbmgGdp/SiA6AP1A70INulGgY2w/ucsGotoo+a9kRXqvX
qfjVNNYSTRJZ1RLPFIvtoQ+t1UoUG7hH1YpmjLFC2zXv65LtpYGPXTMJbw7lk8/u
P5fObMSvux8UUkg+Dl4F9AamIa1uebavbkbhiZojZvJaj0977GIAnrRIzco8Srtn
/UWTDkOjh+i9M4xDmigxwAaWgEXBjMgkN2hIC8/qigCZp7dvem/x2pLBXfngKgs4
dlP/PT4nug1IKql6uLkuDtJqFh+tHo5dQFWmhLJNvuwhfA91X40fGiNzcbdeouGa
3UykSHwf8QfgrYUgfZzSfKCXaEUfkX0GW5x/CBD/bufx74QSV5lRlL2m6pDfjWqo
+XXT8YsvF4HepLYxq3YqU4Fn1MuZnnvO+xv2aFoiM/vg1H0ZErspFvjA72fiJxor
N6XfptMn0TOmAZ9LIlIZdvpM6C780PP+6vsKE8uIKlJeuHfInz9BPZMRyLxACE+T
QVB1YpifdKGv5Hr76mILrNcVQ2H0VuFPFexFRtxSrjxCYXE/6GJXD1saiYpO+EjZ
WhX6toDH243Mg7MzcRdIuJYkEWtdAs5C3zyng5ep9MWIboAjNfCWoNoSTuz8OZvB
fh4lefsNwQBX4WjnGJzWOpEn9WzNQODkDEef3RXBblyCHYORQSy9P68v5Y7AjYHP
9bPOj/CJ6CuCkaMKZq14qFr9YBizLriuIX/r4Vwz3tUHPNDa/El58XDBGLlTRukO
COiMdyDIKTjbwxnEixJoQI3iZqDMte0o295h3hehiVV4A61E92JU41MCCzP+wygy
m10Uyc5Eq0F1Ut04uEg0Cj2tReUCaU2JwPhaOzS7rxZyD10T4qP7CqA9KYluaSyj
RJ4QYbH82+mkgyW0a6UsdibqBLaldcevwYCQa1vqENu5suTjG7OBZzK698kC5FdB
eNT2LDw1FTbQrNX/ShPY63DNBsFF8G9dAlRTO58Tjem8PaIQfYtWTIVj3n7Bxebm
jDg+c5AzS3r4j0Oe2DM5/ojy4MMX0KFvh/NdGYHL+uAyJ4JNH89c3UaHxnmKoY38
r/QL1rVjnc6UmOP+sQC/kZxceqh+FmCebt02UvmhJWOeEP9Pd0tjYFjyHUuAbAFc
HxqAM7/DMxfdIc12F41ndjPxgiOnFatiCwyl6dDKAFAAG+k/Mes9Yfvd0a+L+UVw
xi35uP5/BRnoCZVf1gG+7MuGSarLC2i8v3/npROOc/iLNRG5NB5BcvBbemzK9x1f
wUnni3Ij2edaSf6lMllbS8Zr8Tt7oolCzK5GlT0Gf5hAef/lZOJUL7wUuKvoY8kK
SBcS+VQzsQIsKzGoiHal04nPeY69HzqACYqG6vO5QnohfixjbCPkShXY0VhI0Dbp
xUArAwCdBPnR8TtzrjqDUrvnXUCi/oFjf3eVHDm74whd8GVyPo4uYZmGmTWX/KAS
8xdRAaIVa4T0fLWTPB3TfAUyd3C6v26FG6HLVT6MUNlS4jJNEU9Q4YKT3vrrdCH5
iargL02GvP0bSgwrEl/Rbpgjv9l92oEJLVez4wvFzgrMf095Wq2MHSydqM2/dtSk
HZWWv3BrrKOzX/3n1vfVcbFSPPSpA+Lgaz5GEwoSfXv0YF0579osDcQ0pULNG1ik
vujgDUaPvZ07LqkFQY1YKbmdQmBavhhtNGBS9mcjIs5HUSKDAexmfBd5zuNOnzGw
ftc68UPSMMAjomoVb6f3UJGgqO0EczIWcAt1ILlixEojyeWSvB7ibaCkhd7nbSUf
Ib2pv4ZhuJTFr6/y7l8duyNioR1u5ePCoj1IqNkvBdho0VYmsaxpJ9i2Rx3md9Pt
U/h06XaKmlK2SVIVaiS0JyDSiKIM789mCfGOLL+oXBLpskszeDrbl9P/FX+NXnnj
zHLetqbRtlZXbyb04dataqULlN4pZiczeKex2GrhLdsXHi1Hlvta39OvrrawtVKt
P2tmEuvHIN9OAZBWyvEZcRljsRp++sks6o6obWvXZ3ppe6IWQNxS/UwD2eYaIj5E
kVjf2fITBqHw1fm/lCWO9zQ+804e6nG1M3GASIgR6GRCgWZhjGYwlg66kc3r8DOl
RIRxDDKGnVaVd40XVw2fY4JOfRUqBUqdA1SLJqbyTHYoIzoxymXqId4e/lTqBOME
H7tjP8sPsniuN0AZ30Oi57XBoOJ8Ox4G4p0lrjwszYYFpbbs/IpuInBq/ATEMH8i
fPwo0VQhds/rBVbstmv6ftCXIerz3LKIxnKMyH2TLknBjVtPQxGxXJ84I7CFicK7
GgqossVch1+4fFxh1p3exVNATWCFZnuBhRb1lWPMQaaXaHUo5/FSXQ969p6Wl22D
FxKXbsWCK0vrzq5vRecFlVORUqQhcwV/nYgJwgK52mDjziHfma3iqwAiiawXX889
xgRt5GtZakFJvro/663480yGmhTXjeX3U68zbXffmnLP3wcRJk5Zgg68ILotDzQG
OzLVXlAq1fGNGRvUE9/ebOc21YRsEc5CDKUYPc14z9JsHcWIm8Jq/WXHI1fRPy/x
++aywyV7LKZq/MuEDQ7LGaIp4OT8tJa/5vHSZCZudO3P8qwiCvN7RqJVFopO4OzR
wBl+LTCxQK5++Hfe+2RjKER93dfbu+5mMhVOOq4d+O9P1+4msPM+Jk7jCoKrDLgm
KLx6u5kY0JIthRPk5jkq/YhDUuBW7Vr3xUDx2MZ9gkJNr0RXfzrXEbLjsySlfZz2
QOAY0F7TM61FB4TGKdbSKnoWsSnEjj6fYs/oG4JrmIvLBWUhZG60q2TcReK9Yrh2
zyag/wuXKixJCDeQvyEXQRGDmseAHr2Bp5m6sm9Qs6+nUkXTI8AbN13V0ajKqoc4
pt9HmP6tNE4CiWDz80qeBzzVbUoCh96vLFKaqiPzo1HAq6C6JAi/LEN2yq+uHyYm
e6JtRh50QkQgSA/w5zxmog4ai1PV2gHnGWwjATSkxWyoBgxYd1XtlWTotOHWg9H2
HN5H/TR/sBUgEOZjlRknZ45DyFGCDAXssB/iZ48oHKT9G0WOZRLfDR8L8jvsTcQ/
Umh9lfGaLFf+2vh7SQxa66CsQYi9xOfhrxJQHq6Sz2m9kK2dKkD5sj+9ZBKKOXxr
LTUyZFDU3SPHb+3gU0yVXQf+hLEWsqZyHAmCUNeJsUsx5s7xgFRVZvYSLSL24Ll/
uf/vR9qhV/n/1o1RyEDVtbYA4hxJyfwd7HoPrboQfjJMS7s7OG9t9AjsSv/PNzTT
UaAwumSCevuPqBhwv7KOk7FGonigmB5GYr0PPVNaJnPptQqkeY8QnqnthqZ1f0OZ
MtNV8jpSxKlIhQmsAk2zp/8LQumBOIrX1LZfc66mN1xVGm2XHfC8ySLVkBrpnTYL
+JG+Wj/3Udu7HoDEcTzhhEn5BvCccGBOXlwszAVVAaUVB6p8Vi9H8Rpi0+tNocUx
U6UwIbYLsz7X5WPEGbs5hHdDWmOYHsonoNlrWh3kG1EuggbF9ynSZXVc15OUdG7Y
Srwn+QdZNIACp0GsHQXiNRivWun8cfxV4/F+GwvGJy5oDlxiXAPaYaBEaQL9n1XY
E4eQtFyxy/dq/k95cjzGEoQokGAga1Sd3JBIhYaiy9dKgJkvoAQ8+poBpcroLYYb
ycQFBxWP8woR0k1+NcHWF35Aqc+5a1hYYbdDQ/zzlwM5eAX7/9uKK1dau/VdmMOt
tFtJdR+uQTHv4+AU6u507r+sm1/BRY8YYbaPespnRBUC+UZfN2JeUZHneZ1vpoJG
b6UEej23T+qV2Sh/2JDChdzV4wl5jAaQjn+iH7JbmH/an4xEC7TKheFe0fYuTOJf
dgtp2p18EN5Q813iaiGGtO1y4ZCScKR0hnKzLxXqDZ5Zu2cYhl54htFGhgYMFOJ0
2CLPDMuXoJNAiFucTBmKQVgvGfkwSPmXfhk69TZWuY4iUYHcDFNDVPxInVErDBtw
yiHI0Ua6vh53Ztkw6zhp46czrlZyNZhKwLqZjEXqXCQwWZkYyL9sVImTzHBf6CvT
Z0qmPpFje7SEO/dU/29VQoByBfgSvYRFxaoSSr8O7l8pwcF8JHyMjDj9XfvocWWL
Rg2lhz1vbVGxx1heqI4Jk6RYa78uVQK4+3+Yqv0OHm17rOUw7OR/3uG4Iy9eSULF
kbgyB1Ln09hpRnFDdpmOqEUyi6bUZp21M5+5S108oLaySUFd6ydU6jgOfGYAsl+s
FU4loqwddXexb5np4Frl2b5krEYVIQYPxAlaXN1VnKiF6X9xJo/vnozHTx3+/4uM
erCT66TMhG4nkhsDJpKHmbigU0V4jS/21+WnxP7ZsbKUBCbp473MHJnLOj4XSt6p
pLF3sRPDhk2ZBs44o/unbnOPfCfCNU9hQX/JVw7FW9ffl3gUNittH7q6Pt2DKPpB
eIDFmeecKtEG2ekFnCok63zO4Sk8U/1xrqM4w9/rwK6N0pp0Y0ILIlOFzp3jIs2/
Sj60DJE9tseKegOWdoUn1uFTuRx5tBbzhTGNa8/cLveuW/gFpGlVAD85XVztunGI
/JLgStXGRjOBvldApLWNmEAcdt8+acarm87/ej0BvF5KGghHSTRzBSMVwGDFl/im
E0Fz2of4mXHp46jklmMlq515pkaW6NTyLJqjwM0ScVB/PY0Ps2zVWz81QL/ZeS6s
TomfmAo3XHQxEflGGqy/6owAVmYQHL7+etDlFyUM36TqFofr+mOD9X+vyCTv7vF+
s79qKvKVxzO5UQbGhdjpoy/VLLpf7HYw3fzZZXvj9xqd42hv4hZDKzKvhoShILOt
f2J1mGiFFOr4qSTfgOHDRVNE+YC9Ksu0Mj5lccOnUM3REBXCq7/s1muOh/qJAdUT
KbxIufALPlLvXtC8AsjnSf4ZvSWftTKLEP0sGe19Dm7g6C99Zl5WA6ALpCyfmIbd
mPDNcPMKmqVbVvtVGxmPyI6uGO1EPmPu1NM3woMw0fTqXWDHts3Cl2gWl1UbEXpv
HIFBGIr5TuvkZa9rCUXXe92bgxQpi9uDhpoW5/aSBig5SJCvIw5Fm45Tgy2S40sf
4DwUgMb/TkK4U4CyoGiUyydYKLKyvVlSNjOmdAgJzpnMUPxRucanbahgbeCOlnDz
/ALoGlOgUUhHB5Lqs96wQM/NugLrWAzxFyd9hlEKsiMUWNvNrOUnQhs1shokwZt5
IDkxPqPEIhW9rMqdlkk/Nh7/GuAXAomCvs4/vjrjVV4mjkV2aWS+REMciVgds2cS
G7UYLzjzwBNBUeWpOhaLUjMpDhI/c/CXUHt6iUeOc7u/IG0tI907QB0SXfhvfkcw
J9nIeX6BjnGgJYmSrcy5+RSimIuQpDyUFThv+vNJuXGX2u1lEA4GnnMf4Bdldu+5
uhoqR166GdRwy8uh9D2tqbA+U6xIDEDunibwmKukkG/mWpV9n5vldBtBOnPcA3o8
i6chdqF03P+E0K+oAT5hMrukEOqZxqvUiMmzVX37nlF58BKxVR5NN9DrqjZQ+3bt
dMJive/0XgPvVpRrzPcIEGBO+T56MRXiJm3qnQIBitI12TsGNKQYCyr03/A/dAiI
kLmAm/EogjrfpPvXh8+tOGABJau68EeL0iuz+U3Uxg4eKSC9eT9YZc+zeLyihp0w
kRWQlNY79+RUkzsqeMq15/Vi8gyU8piEROdrEmuRJrLLzjUhficaT9/hN2TElm5r
bYDHuzIowQ8lZnRe1ZugRQdSGZuEXTdvw4PYa5ApVcSwNl3FDtocOy5bwUgETGcB
Qi8iOKSfeznjxn4JodPm75mxdEVoanjr3bUGzr8Yr4kR6znPbxGmakuqhdS5tXBU
djS1HDm8y4R7oWItsRZXnHc4ClW9uQGO8sDL0gMyr33q/8Jl94LVLEDv3TIAuMJp
TrvIctetv6HBO2b6iYKqVwphSSxJ23CrkRYumH66dU+fx3UKJVKcKuQdrpXizmgK
nNVfLDSLQw3Ry86MjIYod008c4zCtEAga1Q2TFd9CJ4g0QsUaaeWbgx9gU3ogIvX
kggHkvFpM4YtejTonOPbJYtQfqBf7G0QNUqTSSgw/B2UrzqgSSgu0LE7MuBVhJ3f
OUg3UEswAbFOSGd+u+uV3Tp2fg2mbMbhn4/+TawcFRKkyC8jsH3sPK8FiCLrbYHI
my79nyUjnF5pBsGLuBz7nw3MNwqiBfU913AnZq2y1DQWzW0NoZmbMijKSxdA2kS6
BS2fPst/QUDaW/x0nyxTc9sleHulW7oVpjjD/Ee05Fj3tCF0N2DX0yhGVuBLyYI6
udHuilikt7HXtDLXHzAb27zZ+P4DZf8P+7zUIZw3pu4fK0GJ3+RDohHUtggRphUw
V6nxMeazO7OFe6z2pzslKGzi9rajnndGZv9reHqBO5jkcr7orqCWuYw4Mwrq+3zh
lCqkWSklO+6GarlOlUaQRFQVGykCzNqZZP5Vy+JkAlwk5zoNmGZDARp7Z+y+IcH8
lrmsQ1Z6uRJm0Du9ICxOp+x8lF8JpGckfU0OYg/PzQkQMgmx+Gm8p0PEO2BR9IkL
R4J0KKSTTszYED6mgDjuenDeao2donMYZ000fBFt5yrJ6oR5XHIGWzTbbutYmpon
tH8uoXvVefn3EfbplkPnBS9btLZc8Tj369/uIpJ3WOAPMEbXFeqf3uUZ+8LSQuEg
O+TWS6XjkYotJWKLSm2jdMuFIpCd/wbbv2IybB7alQtDw7A0uSFm8kWnmfekzLco
HuwzMirSXlSE55yxxWxIbyLFrhp71/ozqZaQsNGBj68dF1WCGVkE8WItiyAT8OEu
OfHXygd9aWUmotvw119VE4F1GZJpaPfcDDdPQuy/AbIydkYlViXmKMi5xZEy9Cyr
tvxOCZaByB1k8orWPdfNfn2bAzpBB2w0kbrSZJ8fY/2QPopo9+yDQqjwOtSKL2uI
J9WJyP1jYoj3CG35EKOGJTui6wDHm1HR9+t7IBsbytn+J7qkDJPLLTqL02XqWl+Q
xnoSoY1Rs9MLp2a4Pcw4QSZ6Gu4aRtlZj3uPWiJh8eroTa18VMXtqzS6kMxJf2B7
NoAsasFBxWdzBWA7fqDcgAkqU700rR1daJSm/+20NnHxggIwFNJl3sTjlo6nkigT
1APzq2QbUGM56zcESl0KAs8bNg7fOLBYzKV3nNiRFhhvfaTm1jARkwLGDdWUHzBk
oPlZfgxyLz4Kl8Bo8EPRzjnyPP63Zgn+gMjy1Or05N1Vo53c1TNYFSVR8aTRUyWs
RCGvaCjyfuOPG8cp63FJIpPzEEmH3Os7tAqX79+KzrgcrL8jQWfUDvybFYk13NUe
MPJ+AZxGfNORnuMQNt+qvkSUFl7+PocI/T64h3WoRjmXF4kMrAKV0hGYTDu8HXMX
NYaJ4Av/ZbjiJx/lAkt0jPueJGc38pSTv8rKVEWZfIURSkYvhuKMcIpqzIxULHbY
4mTgEpKeIZDPcqxcGpGGSdStr9lCHc669VNderJM9JOwJ26uO8UO9B18/jJDP5MB
nVmm1RzYAlaHaoRzlPnTxofDcJThkzkTzTFKRGHVoa8iMXCTUGjpKRna/IZEx/Az
lHTouLqQ2vKcnq9o+eDp/+B5/jaZ+gCxp6FUlLDG8yTjPUXG7HAzsUwnCWPCYGuQ
hpfXOEkVvBIw+/2z7YJVNseXVferQM37b18CMHkdVEORuvMAd6TsHOcx0JVg8Rhf
1tk0zpVaLq0YHhhnqWa7d5ziz1tPrqUhJH+TRZ294ZS0wjMjHFGDU4oAHKdY8n1Y
raMhUKObhyWSAFWuUYmNDU+7eNSOE9DJ++veWjxO1+IIw7ejZYfzh9MgURf1dZAo
5gOHHBX+I7tHnJiIaXz2Osnv8Toz8FPNseo532KYtNp9WJm+pKBpGtdUzDE3fYOR
Um7TXKWRiyinu7okzgcVp0vfgdM2BSIa6QKcSrkC+Hni1V1ZI8/aNWCVzefzg1QR
xiXcivuCsaitxJwcfpH155FNKOFvwx1DveLAN4UmhMGnydUHQ3f5a0sGGwk+i1eV
9XpQem5/gtWjk8QRHZoTTsBpPbRcm8Ki9WEJLO1bXFU+FyEXKAnyhatSpUEnWHSa
eKoyLQzzEo21MvCbVl5tdU4UkGmrHAki+G3PK/751mT6KPUHL2OjMg9UPocXychl
49kwtmX3P0pzPNe4IWKFcInTgFW/jcJ6fjLIvDuxQ1VdGn9nU7YO5KPGsZlQ0Vd6
WvF7gx93DE33HmkPtjjf1be5R7Z5GILMYsLJs6JVJbHeWarvJAK95BO9CbGcFi4M
+mSp+JFWKB+tPgpiI6f0aWUndClNrICKFHpj3DwOUyd8DN8jMQ0gqMk2OZMH69wT
sxRh7IJrmCSfyrqLuPpA56ELIgyVDHOHGyffLuwQt4NdXPO2C7Ohle8aeZcxzNTE
C7d7W5L1vZUoqlyarft7Ru6yqtxBOSrUBsUcDc8YV7FZSru1bMN0T0OnnYuHoJKx
Huka8pRdtS1hnnrErNRLQtNflCgRj6PqGLtIzcbfYHi/PaDIo2/PnHzzxj9bXRVn
G4FtGlazxY3R85U0qVbc8b4Al8Hx+YzmwZfYImu6kC0yI6NLiErOYRZM+3VE/biz
xBEV6VPPeEIALsob9+To3MFZdUwjQNDBV5Kwgx2Olq8GHjEnKIxXaUyD3UJc3sXO
A/NRgf0c1InwIP8MxsDDbx7fmgcnN3O+UPAxdm8Qj46MjcLfV6JMN3tQZRXkyYg4
SQlwq0jf/CGS2JbA5pl/Ebz/cUBPL7SN69ae8u/cVgr1Mmff/IHzUroyF27XXztp
G4RfMLAS4s09TA2YSX1F/r5vdxY/G6YkNv+s5swAbdC56kWPTdWpKpe9tDhdB8hy
n9tHziTA/hB/8ZHH5CBTh/79eu9G/uQ8IKuz6VYYr/REW088crYNvWbxeYljaymX
zz4nE3/BxxnlucbHAO+e1C6SYGh6rmPZa2tbyxbO9smXlnBsbhl95SQAO1pbvQSV
mhRALxvy1lLKI71AKfpjT4owO6kJjJhC1suPGRg87vROCvOApavbOxXzaMDy0duQ
PprSWxucFPyYtuyCCpsC+ArZ2yoKwu65j2emjvFZkfIjjL5gr7WXxugKUEaejAPY
hn/KLQYYcRdm7+Tr5jMpEYT+48La89vrO55AG/I5onvmMLyk0nWBHyo2HGUDYNSK
eBU+Jr4tJkwWFSAEM/WABqF2MtSeGl5PoFygsf7NKRzAaF8wu+8aVAV9KH1qkPQD
LH2Z2/JYzgh2rfQZC0Vllj1gkHK/6nBLjWZdUx5Y7CXczgUhhPrRyNfL42VN+MYV
ynMEauVLxdfslnMyF9D9S94zMCei0QOjlybB5WrcRL59qu5E/P46g1VQs/hw2UGM
dD6dylLadf0vAebMGOsACqIXuVDdewDwVsR/faMgaEh0jVjLUNmqWsxHZOEbYUxa
A7Si1kmf9wXr585I36zVuJAstxJNWs55sRTGkQuqasagXQrq2dvXMNwdS+9N6shM
t3a+vADa0Pmz1lgqjZKeUFcLZ6Az1ahVX9A0aDuXotKyqIqKlue2ADOcQ3fo9R3F
qv/zaXZnnPOjMIDOgzWUTw1Ku7pXEVnXUP5pGkBxl8QZbvfb4NmhZe0nNsWpaIoI
LypnF+StZS1VE71AmCrr6q/TfE+ofUb2P6jK3ChGqaVPWn56f3qRH8B7nkwsjMhO
B6hytn+aYgGnw6neES/mPSBmBvasMEi1+7IEU/2XXpJE++PZ7EMfXh3x1tffjI8k
5TqZu4Jydwyf7t2iYXILPLvusbQrJbFY/qbMslxbU+7RHO0CeqkBW+G2aRUAScN/
9u4uOyV3B1RNbQiZ24opP6exJWgIH6Gsfo97UMz3VMrZYhZxPKufdlXD8A6rhXYP
XaaHXDBeaZUFVctMhkw8qK7doHS6fbReH9FupVdeaRimmvCq7mHCdSZ91WLiNm1t
c/9DOruwD0OwZ7RvMeJu3F1g+oJ91gX75DEix2VeLK8GvWvhoss+fOXss/g8sb13
RVaglwePKpOlpWWxpDbmF0ATu/Ulvwqw4BENmInrIeGU6K4kx3h2tBNTb7lYg6Ve
J/jmMrCknm2X3lGuKzP0MOdWGYPzPmBHWqxYcsQop0e5Hc0/8uZt4OFkrtZCVWSE
LwQ7O0fAiLSUVuhaeND7IoESnrInAPG8TYnPC7aNvhR1YthCQBuPLtz+KUgyt60A
H3hGcgHMW2JQuSWpRa9BeWOuskcSS8V32MykDt+CVL5crbu5pYvaGsliYQJgVcuy
Y4UWdcbLV65vXm0ivdQke25hmfu48c06DTtBkXmHHRsVaoey8d9CTrfjnT59PUUY
AgZtjNrH3iNDm3e6GG4UnHYdwrMr9u3YYs6vKOf1abxSMxT0zzhVdta5gs2vUBzX
45EQGv2HnAJRepuw9da21xe9kyTMZOFTl2OK9KeC00+1j1C0r744iXpHkvLaztWl
g8AZ5UNiRM/E+NcioqmMYotI45htNzGz5oAiaEQxJ8g6axa8qn/+pLi7ATzDC9nR
e/hOxR9aVkA2Qc/I9FbwwUf0pVVXLomFrePeSI1/f40ugCY0tfZYWW6pvR/4yrTo
+PWK4LSxlYuOw6XFzvCBSA1AQLTA50yAsae5HnIkj+kSj5SXiOJIoSooIQ9F4RFf
aABNroOJ9TTOaJ1s0qPss6OeT8xJSIAgSTXrE387sxP+P0tjWEsNTeNvpiUk9kGy
+TgLrs3Zhnm3A4dO+dKvPyiBFhfv2UIpVfaaWpmcOJYVkAMGyoY7RnYGnInnNhuy
MLINUB0eb3WSjxpMBzhJRk0zxCmRbkZcMeISuRwEViuySYmDKbM95NUJQLBnNhyj
PcGKqGk19g3yDBye1Jhf9OqL80EjPin3O3ab22Po6l+fgc8MIyDA11QUD2an4sUe
t4bjzxSyWKtHhFtuCwYfjWPxTGauZzPm2stWaj9uXKowzbDBq1fBHAhz8PYWRZgS
hIXRXhiVAK04zB0dqbEI2RlbVscJe8n6VJd44muf4PRVKmyiC7TzNHek5P8iDaRF
qFkE8FcmBlFzXl44Ptu119xjN8upm/zjcCfe1ISw21eXAocGnhOSyIQsXFpMOXFB
EUge5Oh6XpAR+cvo8Pifz3mPxQLox0p4H+G9dC+VEh64sJcyMdvTvhvbQl/VOrw7
RMEgdpwb9BUUsa50O2Urip5WGpiyE42/fIzyzHKIf7g87WuQe6/PsjOkfvqFGYlQ
4FKL5Jg4+dcf6BivsMx8fyqGYt5bon4qOtiUk3ovyV2jFG4DBiFAMWMw4qUNdkkk
rdjYpzCZyZJxzRWv2txB30CsfgyObCK0pExx4BuSjV5fELU3ojpcubE00x36v0lL
ffA2cIZH1l28VluVKNQbaIv0FF3/zcWrd1tBZEXSKgtd21I1VG4WS4kgaphWfUpH
SOrO2IJhMxYBob8dp2UHn2s6bg86Cmo12JHQ3zXINB8tMGm4rHN8j+Pd0w6pG8UY
1HGZ9478NgxRMVd6LLhgdcO5kRWNbVCJy8bsrXsXQSyff0n+HRyUccTStbUytNcS
2IKPZZDWHZpyxk5CkCK4CUAY/KzNAPyPvi6sCky8Q353/+tNUb41TQabBXiZs1ms
bG47HFgiH7G9EiZoOc3IqOvzVT+0sGniQGRY7bfvrF+Ix8Q5K2zOqC7tZ1x8CQ7e
sI4AKUybwZuTKPWo1t3jhzbVkF83EXVgl8mqmtNFpkHOOsE9C37Ycf60hQTHGJ+8
FCLfNKmhtIlKaF7B/BKRHyjKmap20KqdG4W7bfxTPj7CWeIoxD89lKkZ6u/5bw7v
yEVqkYt5xilrDSA65cdD7M+1cMHDAM/KXlXy2G5dkSSqVl+Zp+kEzqWm7lYDNUEr
ZJVnBGWWy8o7Ifh2V/uibN7ST8a3Phgjb8vaarR36J9cTulL9GeVj+RHloGA5yHq
wwwnjWkTR52K5+IG9MYPrAfdOa93DgcHxeZKRAiTKIp4KXMDCMHm03HMnARt99JE
nQ8rgtRPRZJm/5+3uhdEU4mtjLXdXe8JbcLgeh8gZjPzAaMGt4S//OWwi13Bny9s
H0hekEpm+/WV26BqNdosVN33WUWz6eogOOVlNYdg9hhHNkXZqOR0+XBsmW4GwDmC
I0pZ7MkzSrK08bQr0/EbkExKYdbrfTMIgboef0BjIrcVljZk+QW9H4RROrOnJx64
qJDLs24BpMujNeGwo2D5H0LC8F7mmEU/nZBnZb4l4qBGwnz31BYp7QqyBfTf3t8N
LVf/Wkb6gB/+rqxQakdYEYDA9QAngQK3jpcyH4xLxIckemA46Vphn8EzFmzy918L
wdTOxYA1JBkb1zCFgpnk3QAqlXy/d9yEIgr2KODJaFUOf8QZRPfB1q5/8Zfc7/6P
QBaYvENt1V0S3kj72328dg2JTLsEUCCriFb1ZKsyBLudwV/lU1z21joqVAemfCGT
paDIoV/d2lLQ1ueBLwdu2Wto1lKHQSwigTsG1pn95UaxjdvX86am3lUyeiX7j795
JHsthdjO3m0y20i0XLjpjUHrpDyyMRjjRF2wDvcMRU4H1IRqKVVLQxzYb59LyfjS
oRIkLAeNWOU3Y4b9/OOjZLo8nlIdA6S76nNf6AArdBdz33oQPm/lGTD2nyE6MxoQ
N+0HzIq9B6x0P9n0PQUAqTFeNn1lI19kNjUhLw+St0ES3n4hjgR5IrtM8pGC+kEV
Vh0D4BheYYDPXSCD9g3IA5XNiziqwqKEH9MJvI1EQoCnw87+5RX/auLjvG+NQjGx
XzzQiIziZMOuZ5V7ipCh24M0fb6L2nXGgGfO9Yvw+XEbYC6XyVTXO42B4A5xmXvC
cnb7gK9rp5n/jGmtTgjh59pyx3nLCQ2DYZBIvYKWx0Do+ABTgw7bumf6cObP5iFz
TYeab6yQl5XrW3BQVW0+dB2A9tJSyBVdUnLBSpVafCMuhZKhhtv/hWjdKNhf+aSB
2vc1K31y711+sy1xSC03P/PGxxYLxBAdqbac18RVSqrkYXqzeDu97z9CnfnflpiZ
pW+CUHiLeagTYe2Qt7tVlMzxqcf4pJuV9n96L91L2Y7UH0BnC0qSeETeTzpLPZSP
UplcWaOtgWu6ZqG6Cv9wbPJRSrPuFdTZCpFNXuzZFZfjQHCJYskNgopygOqUtWUF
bNC8CTCmu3TJrWLW9KLtqw+sopMdPzLFgCOWptLhc1HQVi8lzqlbhfj11BcFolXM
Slx6BM9c8L7QsQDSY2o2eEUJLF8LalysnBevFQKhzc5OVfuKOcR/kHiVnTDvJl0g
Af8f9gpHLw5FmDjEvFjt9f8X8VEIpvEfMZbRWBZT1+9WLBwyxd2v72Hs34peq/SG
319QB+shjtQc4eNzmVQF0zmE1Ad5YTrTbAWtm0WONgPWYc6fzvJPSBaEiYy9y0yG
2f9sqtdKplZsp1zZz++64VDOqTEIErt9YlPjG2dLs7TRgFLhj4mw4h6AE3X4VO5t
JBlSL4njRY9XDC11nxq+7cbnUDCohae/uvOJ2aEMjd9fpd4u/sfw9rMjqn95RvvQ
b12s14L1Lo/8Bfq9K7W3bh7FQ7Or7WaAwwLa6OTr0Re+29V12ASV51I5e7tOSXh6
dp1oEcr1BIrxeh9wRgbWTSIBaXz/957hEeXvI6wufEiVv85Z35UPjwEefPfY0x8e
ka48RVKW1YAdwKWzcbv66mOQWmsEibyGgz2i/PsmdaJWxTx4EIe9npwYPve0VLg+
Hprt/n1DEGWbbWmO/irMRSm7WbxDCD5oo2+KyWRmBv7thrahkwZrro2umEXTZh8a
w2YgbD8zK1jF2zQtnWVXJBsJyfQC93DwCtuX8vE8yvztMX7C4CuNjVFF0r5IDq5n
6a/+9z7U8NcneTCuwIiHBOFysiiuaIshVifv7Dc2EFlXGihSmLfTT3HDNWTHHtGD
57RtrcMKa5IZv/nk3afifF9RTFBm/ABjzv0bIuWkd1ZAqh2GmUKogTv1tzJV/dfm
SOv1iBf9ttbSbPDDW9C3Y5BzI182Q3NDXnUiN7RsMGogh0saZfnXERL3qjqHsbk5
paQ73nRakIref8yycPijtWx2Qzwp6qqZZbqL7MR62cMzkVFyOa9CGA2t8o05IAjO
RGRhbgo5DHL5oGvWO7XdttPCUdPOZENg3KjUYvxdAt3YU8nr7WmyPg5nitmCTg3k
w+OSjHcZC/73aWB7/2yN9PFwG/jk8V8LmxVzrzHU0rWVeLkzUKbZEYVHSnRrs/Xy
vxE7e9pzm0qt1tmLTxQTMJsxj3WNWhdx0dLfuz9hvUvZ2CCCXb5k6LquZeEHViTN
kfwIW739jhJUT0+dZSqwbgAQGEtqj22YCImk1dw+CrTDNABSORvTzqJJOKgxS0PT
2Y1j4rsmu95WOSnkKbSKxRhg85JSkqfgo5Omi7chflKg1ZpE7f3Y9D+ymqVWjF9H
76XKK0JTI83hQfL4aKVV3N69Ze37DgHrz5RO3Dud9TWEPM0Lkrq6vY6kK3RiJWVm
Fb+UXtbqaP+avH2Dcd4uKR0i68E3ISsCJW1g+Cg/0FXG4Xk/rfFc3aaRzXeZU6C6
noLCw8k7rsoILAKY9QrfKRpqcwOSETNzhm6SS0rvLpAelEOH3LJQ9FI1+uHdspO+
gyHthOw4M+QxktFiud7VMBTVpjM74mWJhODLEZFyj7IMkIYNevOq2nzuv8PWS6On
EBd5ZkrTLl1v3x2D2WcY5ACjo95o+1avE/3FEyJBNrV/cwBbwh9bF6TAOJO4Jf5k
pF+vK4CF2V9uxsFRHcqqqwiibU3jC9pXiN+g3PpStJBHvl45wk9Be5F1LH4jajw8
SbS8WqbDjthOKG7+gzKKcVDtrhQHNbi3MTgOes+HLOmX1tPkFPo93gP9pMGaKpeM
axuvWQPuQqftcI5CdtlvzGYbLyaZyVtnDYBQZ7rlmD+PPkETlyKqiywBErYmkmMy
TVDiA/sHZ/DFWdTtBAAnSjXpYU6GI5YBdqe5+6t2V4sYdf4cBFsijyiqbkYCUqFV
JFaWMlYEpMFXdDZnlJ2MV9JzeuM8pNGKYZCEai7wjg8zMTJCogRG1QhrZbMRVRJ5
E4MMW4GQYi0J+LmJrgowJiI77a+7fiKiyM0yWOENzwcvdTqBgK53yPCjLqCDpeQd
Dr3llEC0SRlsGDzWwYYRqrg1X1BgiqT8SmJmqOkktWC8T2VBcIqP0GTpiZqob6sJ
SYQHbimohJ+nOLfBbCd+msmNN9wYY4zgMaGKUqpndSAHHfkYK5q7e4zmMAFwNl4S
D83d1tiyawphk7whqTPtymmJ+kdbwhESh3LfzrK9lxAxpkguxTIvCOXYf8MPsx7g
w7P945KAJblOG4bWaxo/sKoin7Av0k1EFTC4iBppeeEP3N067bVNbvlgSlh0jlDi
VLpubrQniz67vnIyFnqeJ7YxTiYyzWylwMyjgQWrRWScTjhwnNKLcMXHQ1I01XYm
zs71FfQvMdpaVoaWKlsZqPpTIpzZygUGGz+Cl92e3wgttYt1JOpHCDfKXNbrjrRX
84iN5kHN4CKYQTu8gXjJXVhIHn6Ar6RXi0JIor4QnzfA16xJqtDgzw0tP9wBsOWC
BRo9zZZD6sUYiSkg1PeO6WAlwjaLJRdyIZbcwlRx/dXqVN/mPFfP1qI1Ysfl4saX
iJEIomef/+NGvWbLlS96LKnFsgyl2GrDYjRlFipFV3rpLbk/H5wXayqHVfaKLY2a
DBZCRChM+YjTQpw/9rU5fGP8YJLnT8ZTBLXhlgvV/d3oYzvQ8FkB3EteiAFkkeSa
yHS9AiQLvC1htzA94rDghZnOJghF02Yal5rnX9/HdJwtMjZ2CBB2ioNSg+RY0oV3
kNN5GKxoE9028CLt2Zvx/VHwk15hCj9CjdhTacIVbc80sOeIhdUR0rChvcEuHI/j
bfmxL8BKfJlPp+KRXeUI8Lh2bKrS1oSSTz+Gu9D3/l5nvSIGmgc7Q1/dBiAfYwhH
EpMPSYAIcJHgTpyMEUem45eEbzre9G5zdSfPWWPTQw44UGQiptKp59CT8kz0UT2L
gC7T/fcFUaj04hoQ/WJ6wDYrMU0AlyS0Pt9bhem03T/AhBtP2hk//YmPU2V7x1FI
orkic5PFVTIUu99q76YmEF7xl9xJkdNb7T/p8lntSxIdm9qzUXNDotQjxbAeBcnN
J4WL5sQMAG8UsZGaktYTdi2zH6kUr45VWRAfueef6vj3EPJOezoQCdihUajOJVat
rArPwUKA81kXN2W6Pzj585x9CGXdllfLqgLhRnTaSA6DPD7CoBXW/84h9EvazC7g
J8UMJulXX8ixiCXrdgMlrNP6IARY7RMbBDlKuC0aF9nfIS+61OAAASe8MSHhAHhn
K9mq95XS9InLVIgNo8w7FD8p2yJ5rq74DZfpQA6B9SkB8K5t7LQ9m0tr97l9rgZG
PvNq646a/tFMcROiF5ssrhl+9r0tGZuhKakfNZA/wsS48SggSBwEaabRr+7ulJVF
uhXkYYMIdR4PYqCkbibpI6Ok8uzETu3o/pR852IrpJ5xKiV1H1iMEn1m9uj8RwzI
ugwGrcFrBwVdkJ994SKpGmHUKGD8XrU1BbrZrjFVtu8HrrvkMFJtwxoL3zqI0tNC
v1OPyr97iJ1LNiR9NFr8f6vB5e9mWG4YilKNX9DSamChi/E7R3f5V9H7JjVSc1XC
8EBPaqedon+mIfK2fanfyv3uZq1Hz80m3lDov+oyk9eMY62bXcu7kt0G1MKyCorH
f1R0sRwdcdpYCbjRkvd1LyW/j9augiGo/2lTTTwxoqAyDrnnStXdS1Uef6ryfiC0
KHtGdMxaflkiS/EzxOv2BCwF5vTUsZ+Crrh5NGvwYHKzesm7AoqRpcbffDizSidH
JTthPKp6j3c0XX8Iw+Jhx0Hzwb0EWFNltYkLYCDfaCm4h0e6zzIfdkHWcDrjNA/B
fSMIrbPkcmq6H7e7sZfmBlN0tWBku9wEI8G1pyHXYmXHzrCXmB7ovD5qtCAMcb91
HQfSZIMViWxKQ0A5zgmrnwltNj/hXqri7c8oIvTezlEfiMAL094IJWtT/ZJn7XL/
k9kqb2+qX/viZnItZ6xQ63dmUWIIYhG6e5E7klUXGyXHBtjUp/47qO+tCHHEIvf/
BL6+GDX8IP3WziSvtT/sUgReG+LCyGEfch/zotFwBOr/4xNbe8J6S6a/eA/w4dKD
jtlfSnJDr1phQ+Sxjv7RuVTy3dw3487GcGfbHUwq/QEHn39fk321iZbklZuzJ0iw
UwRfgBfwM1Gx3n3gK7zDZPQ17j7WQMLHAdeGBOSBTLxiQldtjUu9EhqQgEiRKAAZ
7mB36bd+xkj0VeQGdcrhAKjuXuIcyVsX/KD/45OSF3d6woaalAwAhVkoKWTbcAER
fTII07x2tSf05CiIEWnj38Xtnf+WcaHIz3ovd8rTCPomg8DM0Igj/soHbXzmennI
TBftfqGC8z/d0t5r9DrCaWQb60yM+cnWgap7W+or+0Eo0YFPYLQwglJW3Xfj7UGT
etN4SKdwi7v7TJ/fEJREhYEw1iwCLwCSbsTnAoxXOcQG51h7jjEaXT2qWzf7txvM
J1TFSgNL8dEO8UHzBB1PqQQXxZYMkhxwa8GvQDdaUPX0U8gd/WDygvDg7Yzh9RFs
FqWLAGg4KL7tieD+tcbHbwx358MGvTBAMpErSTOxeOoag0mCXJbBXRGxDjArVcPX
it8ZksTamnwonQqr36kthbZFlCIZOwDxbFVtAh1QsEgUouD1SOMbfA0RvCaQ6ga7
q4tsLbvSl+dQ/qvp1SKiawh1a65J9/GLgS6VsYTXrfU1o271NDt5A3SIvDZ4cPK/
hpJouAPxQIHOJmjTR0f0GoYiQjjlwe0f9khHwunghnW/i+9W29mwJe0u1EgrkEOP
e2JLMehyG8f6fI1pX9+gZemmvYa0BkBSoCh8OY73CbfpL8qiULpljcllqzd3EYdR
yB3VqEYPI6Q09ysRVPW4I/mFvd5ZxKFClGkFLpeXYkiqkI8plSzKIk95V6u9EeWS
pYJAu9igARS3pHg0Xh/8/AbCavpfhrHjW6u6/CGNxNcq2HEc97yudaaSnnTBgl+l
y827B0PwTGXJGBQBorr9fgsBrmTi0e/KKVwhrlc11JaRzS3TGhsCHrmI8WLlpPrk
vwr/d5gfN6IqXYuK7tzUqqJ9M+S0B2b5bXm9JiWG7wfhDV8cX1CNJbybiXkBCVM2
09wcpAHwQ7/E373ozP1JjarpaUqQuMa6oCxlIYsfUPzeD3dCHYwwaZzzAo4WSp14
xICDvQnXsRThsYHQWSSkPT64iBvv8JzistDq/vxqGuFCaSLudXcQFGJOAONOtsBZ
Zv4Yv2yb5aKQRogUd9Au2Pj1Cs0HDw6tVesGqO3Ogyon56WztcQDHFxhhUNo7AmE
MjPmEa/yrJ72wFa9jk4onAi1bqg7ihwbSn41h9Y9RLU79xYf0udwChlgFvEGSYqO
Fr48eHb5uD3LeoIUM8tobrPde5gx5GggsZCOyv2pr3lZePWjazW8BM68X5amEx4U
j4YO8tnC04PqNbdmCTNbsgfVWHfjGI988uPpCEtNiJWJXAgbaa0LHQLfkLHJyWr5
Aer9XMo6C0vG/4jd5fDtZtvJPj/BFacpCQ19AdfJKlW323HthDYnWSXbJhSUim4v
IlzpYpMJ4/AG0JgB4KNjpugz8+jFvMj0hU3Y7VWgkSx0MO+Lp1mN64PvXkTa2OeE
ox86Yv4rcYxAgOxVjyEsoefMkik3AgC9cSej2Qzmt4gpALpAUm3dZaD5lKGJB/B3
S3BYY4CzDxwXK+cUBzOHT5/gqvbEBdshMOa81Uk3mxuzTjN4DDxw0qqvqlo2lTc3
x5LzHg3sVXKXcw2wHSkY7h6ceHbTPKUdX7NQRbVlz1/CN2idfnXuQ44J6tS4A7GV
iUJ7+VuAMsJ0Th6e3x0ao6GY2BJ0Bhib037af51DX6x8wqs74kn8ufIqanupb8TD
3DRlWO0iA9pEsvKMlyPJCCSONW5zUSpCi1I5qOL5QDuRx/aXsFP+HBgt9oALeAbT
ot0Bw83SKnAM6SIdxXNp286D+g3ZxC9rcqx+UF0JphsOxFFTcLEIDgKsce5zm3o8
9jZk8LhST5TK2RnwmVj1BmbrPw/eEhynLXcP3XhnDIidVIKMEN99qWL0UY7Lq45g
P8QawYQrtf1jL+kbIdMOECOSmi2lA5fg4PQ9ia/03kUe7AMqUN6ymU4OE3PIJJmT
CuZH3yIdTQT8z76Canx+wVz6eM7P6YBdYww3fpayV8QIDLvrQekIqO2sXMCfxb8W
ftPrRsBKS/URBRUQkYIYF7XknoAI3+67t7ijKe3aryL/9l0m+X+d4/ofQyUa95Lb
N5fu9VQXXSki3UtvOsIF6C2XPkpdpgv3si75ycgHDin3blh0jykSdyhx2qrmRbvs
PuP3jDPSBvt9V90tdD9X9u6EV0r5TxBQWLxIJnxqpXnTR4brIBWtub/WYwXMKZkk
/1NtaGL7yY4QRg/M1jc1jLUnWylqalvhLhu6ZQAF+Lq1MYfSE5e5PQl60laVUNl/
0O/vwzUbDZbJ0D/hK5DD9zFbWj8Zb9HGT5GTogDSX88TvV9AsABAr1MR4IRG5eJ+
2kxXy+9Lc0bQN52uVzLSVGyjIlz+vrXXcZhip/snQC8P12m3ppuvUz1it10SYaTH
WDQdU+PNu7IerdV8J1ZbJ92Nn+BVbz5wCBpstsY0pZcDgiocLo0oQQnKlBivNLgC
M1vIW9PuoqJn6VNNTaOZbojJBViydy6oSoUzx9kofbEcStZgseUer9EPehjOy+N1
c3nDpu1hQWV7d9AyFrXN9zoxKdP2PXPg5ZZhTZD2cwPbZXJ6r8KxHkJgCIMhJE5Y
LcoJJvceS/P7wmX79IiVYEjb17D+ggFhJ8XwBNmX2AE6grlB2MhzeBgQQbz5oA+U
qaTKv9vVTOzuIAZgH56l/uWIRziAoys0bmh1uw29v9lJie7y8OpFcfLzuq3keygc
gD87lLDVWy1F0EsqKVOksQlqMo5/cqu+ysb9v46/5rJf5/lI7e4sUDGp5XuCpvTv
Zq9BKArVfJGmyrGy9ldqQnpDxl/O1bHUQ5a+YrTUY3O8f/yH1QOLBhGO1H5SqDyj
7JtMfcnvgg9INspAghUcHGTa7hcwbfYGAD/AuZ7a0KWBIstTtoryJqF7jVdaugwl
QQLcgHeotpzmNte1950xBjhWv7xZKDlLdMUyW4UMV6QYw8esBlm3WuA6CtBwb9Q1
i3J5nVorrkyfbt8kvMjGYrf/tW2iYlM2hRXjC4f9fXs7v5+9SWt/BZd2lLjA2mOW
v+LkqKQiWdTwbJu+8lmF5DyOe1MsPHKX/8jSknpEotFhn9bo++ybkuI29HaSJLbx
2n/rXsj6gco6xMkrsOw4mawppkHfe6QNlwaCoOCfekIstSep1wkAgrRjsb3JGcRC
DOAPvYBE/bOIiW6HoG/F3kBtsmKEYbMR7nyRHYa9+ADdIm1X8QhP7lvCbbcwQBgR
w5wjmk2R3whLkicyjJIJIqat4OA1ByfwN7FvijQF9B5eSqyO7bmXj3wfUggK/6U8
8Jy0QFwULs01QfXKgoxgpGpncZlM37+fGcwhy9yNNyVEr0qJ/JVaOfZoSs63VKdc
2PoNMrV7sPyFLYXSbwfTaBtlTzC270yopMRT5rxp0ayVXY+CIs3s3DplOb4N3N4f
qbAOwSa7VrMXN/1p6PjZU8AM15pK4PIr1Aa3VLjVudperi0Ti4U02B/DHbufjT40
AVs+4TZH8I5+Uw1spf6fXIoaY7XFGYPx3rl233f77t/DOYhujlI0xwv+g6XL3LIk
8hZOxEgU24cOS8iPv6ds+emDWBCIr2hJwbILLEDmVnEyEbRkfSQvL8eMnDfpwfeK
1IwJH2ZEGSS18QwUGxOutxWrAdyVifLvZnqgSu6+TLjZxB2dqDaGW5GgxbEV/c7T
XAurkdsk0xcNW2NmSqtu5zsPZualwtzNPKVNLwa2hcn0xpvfK2u2usJqej4XCuwF
E0Od7G3I5Dbgaa3mcjS111ADmBN34W9SpfOnWsqZHDKmVisDEHQEZm1eLCMCSPzL
rue92Q3p2iG5x7JRDIMln+w4u94cug63VOQ9XzUN2kJ8+8TokRQG5hBTSX8/HTNd
Qr+fo8pLNFEpRU3qBa0xsTrY2/KI1+mWcfh1/CxViSNdll8qGzFvY4OzhYpiqbuo
ZHt8pUmo7H8mOiMk77raW82mLYVEDjCTUxg/J0T12+3BgBXeQucduPke/ch7p40w
w6Jzc9513K+ViU/pUA2xDUgu64LTRTM5t+a9RDox9iaQ2rD7vTT5e9leduHx1rk3
2VKlNiex3fFU3wNz9I2yAHvYA/0+yRTHA+OiDipKFyaiyCZ9sNhU/av2k+6d0R4H
bnR76DvT9ndWOvyTMlSYLFj+WDGOTE8phbIb6N6jVprfYFE8uQAkP9T9TX0Ou8cm
FxWiDUTtJtyzML9qoRQvTx7KMRqnacR6599QbGqV/qzAiWBxuBSVBRW1wO7N0IB1
Ta4xTckaq1YuEwp+I4tXzE2estby6O+pnugE2S/487eEmQ8a+QDx6TW7Q9dkXwqx
a+oh5z0+zIiHHMrjznKLUc+Uw+r1N9UJHG2RLFbd13COhXQnZsv5ulgTlYiOET6T
MFICSkT54BamELzxwdLlBykuzAVvujTlMex4mUNYV5S1WdrRczo/AvGBT+H7cXpa
CM7yJAABmpYf1Tk3OW2oewOspQR3++RPRLOLIZkYCHnG5ZSOCst5OjJVQYJ9FIYD
MzcKnUhliK/3WJYRpqoAVNWU9lHBl+ANOmbsDFvHy4sbxS0MwLMKRzlepT8r0y1P
WVnz1N4GAIs0l45TobHWVYZU33+LWLuvlaDJ+crpCbVzpTtVSIw37YxAFWvV947r
21HEorqtWKSeJhxWKDUyERFw6bp6jCP28i/C3bu3jxSlYqzFHohq1nsgnTxAMDL+
jWSJ1Rv68kObMT5b577onJMY9lw6MtAc4SpKoLZLs3RSgmvjwSgciCcD/kcIZ8aD
J9IILxqh5KrvJkOR3GLfOb0gHVj0t8+RNuVmDeUggaJRVkAc+62tCCfbMjjUDUvb
D0ESic+v1V4e6nb/jzyJ/bzEWvLjSdycDC/t5oKZB640Pz/+R1DtPn8NqzZmx/u2
MtRaj+1KF/OQ9lZAOIzIRry7+6VcMAXyC1uT14QfaXkFRNjmAjyGT13ShwsP/AHD
6tBHzpalVV3j3RbSUWXc0IsVkxKNo+lHgX1rwYbJDqLv1taJqXyQewzZyIthUcyy
NiDLFoAlcqoqvFhvoU53VmxJrf844X4zMjSnVk3mQgAD6TLQ45WN7xGlvb2BIRqG
g8df1QxzHzM9kIO1aBukXiCdl8vLGaiDU4da9VW2DolYBpe1JzMJK/HOLTuvmJNZ
m3W41UcOoe8ONOkFP8bGBTxNRczOEjLcAdZPGZT6N79LxdYGpmMwKCizX0N9hbAF
SX+ScOj6VUTOmlEoSNEz5eKoRl6f7L7o9TCoGet0HiGguYLP31wrD5ffXy3bW/rW
ZyzWE5d4pchbm6PZNtG+NDoffnu5EFFt9yQJHNmAO9a5HvIMuzWFdDo1ad0vbCMK
Xe8STWZyNqhWWFOsZjHswzhdO8p87O5CeuuHNUc6+dw7JE/NOINPWpg648CrZOaN
+SLcfnI6LEJvBc5X3PCdZHK69nB/80fquVMocEBs3sca13GL6JKj1nJtsNpPOnDA
dBN+pp01BpIkA8V3vpuEhdxCoaTmtDgvQunFhBkpDTv3hJKsTRYDz4hqlsHLFRDI
ufz7BdC3OrLk++ldvJ0SwBZ5oj6zVqSQjqO/B3IlBf31JduddbF/ZiPgAFZVqGnR
Nqyw44GBEzw91dt5TR2RmfMr/XX7qPlKniBJ8wI5QuLrG4w3mDT9QOdaZxo8vP8+
iJCua+tkB3EQ8smgajSzpK4BnnGFqF3UK/lY5QlitBQyZ952GU+ClZoHiIOH16Go
ZvxjdiO7KdhDP0x+TbE04X7thSbDqHjQs6x7edN0rO/kxlinxZiZrBFSU/jLWiry
MNpQsRD6oWDW0suZ7Z5vYEAK1zOcjGDdRi+r+fDSFuMqCLzmPcHpk+ERen83TgCh
ySS2LFeiYk28U1h5/SVgtfwom0PY76xgAehkN2zRJrXMFI6rtA99jUMsFCypHVqY
RlauvadZOBNLg/OXdZQQBBkbQEggt7WEnV+oD850vzt7cRT0Eq0KWGCQ+K2lJoTN
Z6h+ikCh7LfROgnCvmC9JojbCcsHO3aP2RqvZiNOpz7THaSYskbCY/z8khDKlsr5
jF8aUL3HYNz58SpaXmV5Ike7ZWG+i8qfNER6LDTDYuPgItEt2fM9ZKxy5W0npnT3
/ZpeNnNHfSxJz5zZL0YU14C4i1NTT2E9IEGM+otc8oyWCTyevnHS49aEr7pHYrFf
qPp/BRJN0yjrIJUAtrMr7F0pQullYiOjybC7EmjmX7cKeU47ag0E0zZAod4tSjkz
Yau5tNZxV2puw1XE8cZQG8o3dYpSXSuLHJh71Fhm3MyYQdYM1qWU2Fn9ZeIUJ8OR
Zdh4e2St+29onHBCNFDvCZOqS3MieKVozVsuKAmt2PhZpyI69UCFS2VP2BbyEKfc
YzzEWIaPaquSyJ1nJgNx6thIZ4/kN9SDhnsC27opycip/W43i6xsqc2lwM08Qkfw
YB1weWCt3aSKUD9Ng3xpyX0iOtxw7Og/d9KXA2M3zNlYGL7am4c/lW7sM4cpf7hg
tUUoAHqQlngImbKk2UMU3q7tD6aClvYxIJsOJ5F08DwhQc5Tg9aM6cis1bpNZTv/
E99x/8Hh16o8osSgshOROi824HAjey+sjZl9r9029XW0yxNCIUpfScP1ofGlXAn4
NneD8sWlOvDoeH0TrzbGUCf6kopBstmAlp+gpO2HSl8CXexZ3NZrPJ1j5btCeuI/
vlQOibPseCLiksnEHTLP54O2I91VSYq8c9pYdgCDqoTMV44FWJfw8wd4ReDN7VDp
ClJOchBzSAozFydnfDLs+l3+M4RO5sMQviF4QWwCYksjY4EAH+auO0rhfzz8DU3w
A7y/sRT9MZA/KQw10MIty0R3HoGKnQly/Lm17Y+p8x0OGZ6DJmg0W9wQinfprtHS
vhCp5g1WZgdsdO8GoIvMip+JVz+ORhj1Qu0fpUPI/AIlvlSVXG8nA3yYx9P9iG5k
G0KAAxL8KRlwVuD97rzM5ZTdonM2/t6B/DveeFzxAPIMCHADfv4d185fbyAm/1Tz
gCJATHgF8+pLJ+b0uuKvBrvjnAB+3HsJRDSO6ocfPo0ipSqAUtxi1RAg0Q719ecu
TnqBj3aaoL+mvo7H1m1xQWOKjUFlAYywX+aDdLJ+biEycEUowzJVy1oT13OUI7Lt
21YigVJAa/r2XnGW0pUCRl+b6Cy8YQl5O3PdmSGmmACpVbOPgqSwYuDjxFpyX452
4l27/CdYI6RTdl/FXAEsNcM01CdwEDKlQxlKDkkTKTMnLFiW1of5QP+IjfPwLBeb
LWCNnbJ4skgReF2cypc2C8q96UxNFcTnpXpcxvFv5oqEfDLSfJ10Qq1qUb2JdIk8
nAHAEi/nf/H0nJiLes3WEXE3qsIVoiD8a6C83NTNG0/MzR0wuXP0gUfeBadzeCAC
RGkLExPAVOICgGqOJ3ULlMfu3GODgOoQ4on9bsST2eqASV1ukvrY5K2iyP38XKll
Y/1Sv0P0OnpAkP5vTq3cxzUzJgVtCXNSN6v7ubgYK+eEgoJHghrh+auVt4RpgvOo
2bxf+pBTSZ3T/Cv0kF5qlXp+KNYThqWmpD/gCpYZqv2apCF7pNBWNUJVutGQb8Sm
NaExX1eDBjrzJokh04Wp7JZrNy3A7zfLI34zq+NDfQ3+9FwdoEh+i3aYKLay+kUQ
k043L6vwWs0+VAmzq9DE0xsSK86eTpwhpi3NptOv7KH1gBh8KQ5i4pD/ki7tzwOj
Rob/Nc25aUVGSMkuPm8Dzdm6Rai7z9owVP9k+HAqLKkIPmc4FWdlYEj9izHSML+b
4T4/WfnvuRPsuP+8LhppFZ9VdJzRYYly/bbzLpa+MGJftlZ+TajeFBm55oYLQiLW
ttwCVJoyrO4LYIommZODIUP23fgRLQq471OFHZwpiS5KqqYlTJxamMnzWqyby7xJ
l5HwD1AhOZf6e8X4KdAOWdHIbeR+Y9BEiCjGAbmb1hE5d6o4hQowSgmVQjIgdNKm
1LykWojcb/aPcact+Tb4BtrEKkDcZ8iYK2tBBms/fZqWYKbyzeOCZcFkgD24D9Wf
v/HJkiksucQ/gf8Um4hBGSUgZKt47hQv6xBkuoP5Jy2jB5Ia0Y/WmeJwvzmPO7sR
8EO6hogzytEyTKkcFOHIFLtmOz1QM8cYxuV1rWiRvGa7eL17TCdeGG0qsKHoCayj
WdqR3FSdOMXo2/SBrv//YrdH0Fpe4RfvEDcuJur3AG8JM/IcsbqJzJF1V2zKUXxL
3C0oHzCO82021u5TnN+80TlGt2f+Wtrcgajx6nhpbC6nLYrOiTIhD/iZ6S4G1S5H
u/VHKTgoam+ijY+FL+8Een338zPVFuPwAioRhDhzWrJS7ONFVL8+jZvFMmIV+1f5
3icRkuI4TlvxzGzTDayyQbexN3t+6KNbdiE6arzHDlwTCFsHojskgr6ae94ZKrhC
gIkSZQEnDQWdw5ayX0YxMpY6j6Plwdn98llQWLOhI/7NOrWLMXeTlZ8+sYc2B9Dg
bOObj3RMyimji38OTKEjiBnGNTlyf5KOUAOOQBnS6+TRHXgwtcERLibJy/WUFyNq
0Kl4Li94O84CmhcTjK29XUJCnfnWorkjZOzlnTydrnQRM83+HZTGvrX+RlUZE3qR
yclPodlvlMASMwGkcTjZulpG9KWp/ddHbWTKT8mG7lkksQdHCxs7/2XwKiNKTvqv
Q86ZtCvaURFmeWrNuRqrJ8KlRM1b1xTmHw1J8xy3YUbAj74hPfyNGSZvs/rihc+8
Lh9Fn13R2POeLKGCvDic374q7iFgkz0wHlXOz9PKdtQ1QwZOxz+Kjc/pym94ZXZU
u8nGpIumRHi7PiOb5Z8Qqvq5FUMsCe7JZwE5SW9PBhDozy0d4BHDv6EZBWZcJ+Se
KKC47l3YhANzN1n327tpLy2dGd5aFbJKeGAelpAmGpg5oTPKrP32VzDLhdwyHusj
c2pjw0vTxBPcKLkoz4hiTpoH5OmDjEo0h1X4gxPbIn4CqNlJYLqsx4SAmokco5gg
6bMVopH89+u15hkgnlCrPcd/FxsYHKTHjIlbyZmJqzpWjwCf1ly2VCZVTeB8a6RP
54Pes0RyGMOj0x6W5busUru20Bc2r4bFA9DWoAs2uzmf8bfATaaWAnLYXcCt5eS6
LfpV2j5WDPD8lJ2+XnMW39pEImBnXZeco7gW3HtwZiZA7UWOZx/GqMlNwMxLl/sk
Si0hX94I8fQDnSdsyV0M776UDb1frEe2vNXlxURzikwv0mGbsfva/pAt0AFREZnV
u5vOULbTuGbn+yP8mipBeFo5PnnKaaRKMWvzPZ5KrbuZ4+dV6SKdYuOPIhYWHwnG
RzKGswAB4hq5Gw3m+QNJ0E+wwwPtpofkZ66dlBZNGC1xoE64dmMWZ7AS+Llqf8Lx
M9gmYng01Xs45YdgDm97iYSi4wqM8dXRVluFty9S1RQEqrX70WpoXgNV9apJiXRK
r/Ku+qgQaRMNAbzszGwxR/zRrGoZNwNnKrL30qp/bAFHYnJd0chY6ZFZo2he8de1
/9ZKfqmml7w0RrnvmLUHtUnIiQ8M/IgF4QbTMmYSZtDyWXXCz07mSuIW/oYbIS/S
95L8iYQfYhk92/niwPtHY5I0wwqDVMYhQ/CeKTn/WPRvQ3j2kes1GLU4xqxXW5/P
9yl9cM7/H3/xXJ79DZb8k+EhdbNm6xCMa83ZalAjL3/F/br7DdStq7q6b91MduIp
VI5UqgvObgJ/TWj/l0NRO2liRYuA0bcbA8ua9munX/j+rFpZ4glB3jI1q6zcx8Bv
ECMbNAUIOA4GDJ4UTVH5Q+OxIy8uxF2glMawkkG7JkfpzaLECxLCXdcZkPrTS8Of
5DSVV0t2NWV+W3bt0X9i5KFbXSkqcFqutmpEpsS7dfpkMmd7oz0PJSRPsBlqg880
QrNZuOlaQYv4AyqsDCoPIair3PcjOjPv9WSaRRba50rF0jd8YGo9qxp3fUq6OEhQ
hZTnuCjgYjya2UcVHsfVcr9Zl0bgWGdeBNamtu/XweQmgyE30jTIJN4KHMRtGAxU
yuisuNgC/au5NVk2f7XOrleVRB5o9W0w59KFCTSqgfkoFs5UZzOeQyXmvVLy/qvI
DClj59y4gsHXsgPUuY69Qb7tc3CZg6QS/4wk7/HAZPHB/AfWSp7eMK1fdWtVfYPn
WTGc0HXXVrbBDjOhK1r/l4UKSc9sJmwb653IG3ptgeidl/7fk0+RmvYt0CjGvehj
6jbdiQI11DnSG3SG1T9OKkhJy3QLp+cP8tZuSoQHwUKhMpk+XbJcAx/FyDfncIX3
V83sjY0x4USXJ9IjZe+muk4Z4zTOLdgATJh53iYbH+jkesC0eShx/ij5p8wiJqep
truo/SyLwkXBCgo9iqwSn8rlhzJf3JIMCDUekccKbvcdyEHAQW4ZXBLaYxlnjE4Q
YK2TgyerJa2ReR3p2Fbp4P8Ebf6LSPFE2/S5fEokvfwuw7/AwudM+EDAvzX3OYzJ
wSwKa8KVL8vcSmg/SL7u5+5R4AKiUJce2AG7LOF/JcvI3D3F3ljbQNBrIg0J+d1F
HYagC00O70qxe/gw2TO1jQarcSMnBH7/iNu1bmd1qcBqUIgFYY8BFcxVGkd3KrdE
8uiVcAvIi6S6BlfFSQZP+PAp3rQT/Iw80yniLP2o3132nYZevsMPLzpK91Am6Chz
cyZ7GjxHSWzyosa51e2ZZHGCkqo9ArXMlKViCdfFl42AZdldGhIdsIaoX+9x7OnK
2xsd77Et7XjPGp79hQYPd6ULKQMq8Urrkor2eGMcUbfqzfZmPvAFaGaJNjL00far
3nzwBWmvPfqMpJwqPP3JwpGUXjdy0DIwImanuDMRcQpKCkErRLwGLvQAzZy2ILX0
0+PhQiDhLjjZpOy5oPqS3Pzvd+VQaEs1gb9BXYk6S82arRI2fII4kneytFC2cp8Z
/g5TaJNSBQGg+I2LsY5+hihDSdNuVejxK7dtkTHEgsptv9fq0GOGUlcXA5FPI0Hl
AGWhM6n/DmzDMgxRv7mI9xDEako/fOD7+mH/jtdDY1UJVicgAqzOZBtg8vDpQAD1
sXr4FlIkl9Z9DEeX7t50Z7LOpmTzCcFhhD2uBfm3aOe0hA3YQtAiB60HEVWvUNHF
MLUG0KlmlFbePDvJEhmIgQuEBBZuwNnuQWtBcDv3HKGwNXBIHZ93hWXrgEZyf5Lx
y12prsRPQadV5zH3I+eVD4tHrlBhSABBp/lO9ev/lrgLXFr5oSmt1ByvqJvP2RxX
QvQszfiqBF2L1FR4i7jdVxf2exyC1K+RE8BxkW6E/1I8FqJWlw+YEw7+Ky6vKUf/
J2ETzRElt/YK9+n/8D309V4mB6GIZ5nAMJ8dJQtiboSPGfPq8xHRQwXKi8DAKNr5
c7+CWMkbBdTUktXcjWyCM8axO6uZmPuEed5VDzmTUjsWFZP7jGQdB0GLdEbtLR+U
RGn9mM4uq0SyBPopP+OVibN8skBCsCmrhmWsG2lv05tb9QJew2vHKfd8NQXVfVPd
pQ7wiiD5yYQWUAv+xafkgAPMwSQbyJ1rSHT0gS7xKYJjMzSmjwbFzzKx05cQqU8o
0zbLkfT0VytaizGXTl8zluPXTnV/W19VkCIyQeWZBhw35PC3T6B0fHvMfAqlnKeM
iPyYTgLKk54wOeh2FEHcibyAbp7xWgfZ5fmZs85rmqmhW0b/fAbwttUS5Qpkk21E
ORLJeKoz3bN21fbly5N/xnxXFb/zEtnlGtvDlxrWesH7o108wfx2gdrCPjS4kNuf
qOfrNkFabMBWxklJDNAxlDOqnKVlrIpkgOB0oOGXHw8GQcSeeBGmNNlod65g9dhC
UG3hXT26BjtL6X+9I4TjD8P109f7mkLvdeu7ThHS21VeibWisjfb29yey/mXBDVQ
WcbWPT6+LIss5RZY5CBPbwM2ZcTq8FyU7p2Mz6405dw8LDU/fafEXG/uhV9Pkg5Y
n5eesCp6UQSe6ALdZzC/fFdp3zvTEGYCU/3zeCcFefy+pK8cXYXY+GDg0gmT49RX
uUwDOVyH1hyvXA3+edn5OKyWL/DNfZ4p1NxTkH4krucHi7sj5AL6qMMiGBds0+AO
8u/22aPbkIQnlk4NxZGhdrvTzc0TjhHCD3jzGgT/OuMVTdGRwFzPoNeCsG47+ZUy
hz5tssfTGfMg6FxSadMj9Lz3dhOTrK2nyRY9XmrzL+WGNMfSpy+TcaYMeo9fhANv
YaUAP/ktC3qKpf0LhVxVahs7PBPOae0WXEQE4MXJs97FCzmA+XkDpu0NBsihlwsH
rsepeJGBUPxUyfVB4trU1q5LxUYMgJ0Rs1gJwGZklt/PE7XvaAA+3HHh6c7ipDL6
DKHsbwp0mHqKcNyHTYP1XDTFwrt+bwQBOBrZtcVwa2u3kb2iHwFS0QEBqR9cSfMM
0cS9AGFjgV855sddXIF530m+b1oDTqTk2bVNV/9tH4SglT+JuCHQtAeEMSZYTYwt
aU41xkyZ9U0xWQQ88MjGfjILOx7UI5FnoC2s47W+OA8IMQ4nw5aY46AinNRJIjR9
63TFmX37s/OQo0Sz6SViHqupVZN/+wdamBzXkc2AWRNbkUO+Y+ACkxlJsjwezRn6
cplK3xbRXpGwqHvMe/oJy65cGoWbmlYgCaja7HmRRY2rUr+oaku/fce/zabHNugI
Txy5Vk2mvGWZM81LF4ia/XqwM7sJm4pcNuyOJRynbBKvOfbVtu/ztGRnNpZMtAm6
XJmkQn432yAZLwWbMpxcLT3MtyQq6cepBUbJKPePFNs7D9Z/r72AYqlsj6ebEZ3P
9F3cl9tNOFm/WaLL0oQ998VPCPprjzKZPw5bWrDZc4AW6xSVyXvTFjsHA8T8/dtT
FJV/ejByzQCCt/rlAkkzrzP9B85cseNmFn1iBs6LJh5gjnMlbClauSDgUblmHO4T
tzFGXbqiatXtYjC/0iFwc+LLanfNFmF9xoj7nhxXE5FNUj1qkiXx+VG+RBFc3AS9
A8w6U5JsOD+SAFx6WEEd9cHmjzGlP8/055Vmrdr1xFmWRvcUH0uE8GrNpyraagTS
zEg4oL03GEcBnZZ4eH9DVbOYAK3kBntWlJyUtwbrBgeEy2hIjqoGhJCu5CT0FJ6t
eKz3+LSjcYIoqYwR5OLuPcrfjTK+XYIgYbXD847mYKFRjfsiYUYzw1hQmQ7FIp+V
gZrKz5Www2TcmSQm6Xigk0lcCS0KvfoQz2bNDLb9iC8g1qVgrj0SMwsOChiKdpQH
oxc4qtoxw0C6fSjUnvbDsl0zSQwzGcsi4+xas8k9xk8ys85WkcRJfx2AMsCvJ7Sv
3ulq7IQjQHB6LdVbatZExF/8/9gbgDcubC+mb5i9tGMApfCzvD1FwXYvT4VxKviX
JbxxunULh4U/XoXrU219/NQWQNa0anLAMDvXiyE8+ZszcTlN/QWS9nZTACOOHxVn
2g5a257rdboikQcwgYoH0Hyv8j8JqAzAAXnNdEE8uSw3BzreFgbbdwCCdcaiIx5x
I6bEUQKgroN+WFqYiEx1zeVmL/oPIcI7EZJdxQaJ4jzoc1gDsz+9SP1MGLf/Vl5e
jgPaiaIbnRR/HgtSAFLfhVOWO2DsoGA/rCVWzceuAHEmWIMSA1vd0UvuYmMLPV2Y
9bK6EG86vA9gNlDafpipqJlBg4re9PwzPolesnaaDa7kjK0t8zq8Pep5vRjxzFhG
5jhsY9UxkLNKAO5pJ33dAFfLPDxWsEgiaM2+tHvMm3AUOGKjsVvLt7wrRvRcrAvQ
V0pk5FO+nplGWJhlyi8ShuQDTp5IT4QxIzVP9NdNUo7DGZ99KMr8kHazPgGC0Xxx
Dj+LFsFozZafwylD2w3yRmHeq2xQu9/W6U31DDcWUMaR2XYUILjgHEyBK3W5aM1x
s9Zg37n/ULlfg87lUdCWXhR7iqTtS8pniV6sHI+kcXwIM1svpz4mZdrcgM8VYwok
CLZUK+ehBTJrAmTUTS6sRHvq2erCSD3bbY8jgp2V5InwTlOAIt8dY7rV4eYsVDGk
FzMgRQxMIhpeWig4L3O/Ksz4PVLSiAdEX5jNmeAJr3MCd1ltW1wWxnO9j+2cyr4c
0NElvaNBWpqGuRxgYpxCmOgxBFnJ5weC3eK8SP8kfXYad3QharyLkWpgqJyZbs5Y
pfjzPIdjE+biLD3t4oqd6QHRNe+ZFnYMZ8ouNpcwL85HvYrWLFW1LPJKVx53ALMN
ayCe21Yp4MY0T513ka1HR+AKZAMeNdsT9TDAF4SKS6asHs/iKtL2GgyuazYoe3n6
4dZjIEjsSKs5qTmh7jBvysQvU+ne9Cb9d7RcHwvYvqF8C1p9tUcolDNj/pWH5wwZ
clZ665YqjhUW4Kat3uHzcpfR4X8Z89Pa3ec4ulGvHcMV7+2Leb2bCh11N7kfwe0v
lMMv2YOUxeQtuXGXDNfQvZ2RVhTC51JiY52d1TPTyXJbOTkxab5dpgW/Nt+iNA15
8LPYofxaLkQu3FdvqbtbhjPUWGC72uLHzpVFtVmYB49IWd0g5F42thBUmuvsBiiu
qIILF4mhZ0ZB34+73Mdva7Wm16z/oSSDKPPjjwGJokHMlTRJalh75VzjV2grim5S
9junT+DL2DP5EcZivb5owABJrRH906VNlQkEDHxi1tUGfEXv07NKhlLFIvME0Uwf
PRReF7AY/mOpnwHSZxnQnz1ldm4FtRZeVjYO81hTw7xoGh++cKZR/kDLluqJMCWs
zOSZuT/KXB9BIwiVhc62GTQCRxU0D6gHn8udGqXaQ3U0kL6Et5Nm8JNUxpU1T8rJ
e8BU8Ls7vRCrlLeHZodQWjA8KrKmFZre/63mK0xTXQZJVp9s2mLTCgDf1nn3wzV5
N5IlP7sxbzYcr20chuq4CQy/kJoM7+zdAOz5OG5BqZgNl8tjPmb01ZnxCQszlGzI
6NISHEIQ/3dve+6eceHkdcwnIcSElYHipGM/B57+N3QNOhvLBFX7i22icPPfaHKx
Cwe6FvHnY5wr/2wUZWSg7keGvWCogbFaEsTHdhJHPmFhC31NWTro1AgjgfaTceIN
jqpWactiTUuYZWfAMyeX4xy7b1pX/lXU1IzDx+IQMg4mdb7CV2hjoA4Q4a43M+dY
jW3uF04H3c7ec+YWI+28PotrY46Wd7DXz1JojNejahN4pA1uUK1Vg7J6fvcAj9PF
YMyIPDniKkdNEjAWEFNIM4MJeVk5nHkU5kPRtC0ycwNqDJC9ROBkRTGAUmztaGgp
y5KKi5VdXzS+eO2SmeP++aWwnzfmvzBuGKhZHAvA/ycp9zkw/+PLvDtG6vl+oTUz
vkTX+dKrFb7wsAlMUNm0ELTw4SUJY2j7SxMMWIwqTu7krQsyfidjJZJEu/vRIU3g
IbxsY3olLdLfZOSoovPep661bBosdRnGOHWLVlYtsrnFSrUpmQogH5ogPdOwhbH0
8c6sq+OuB7S+W+tOiyrbs0JORtgfNjx7XRaxOk6RsQFiAtilia/91tdm1ibDHvul
OwZaiaA+I6xwqkjZDCN3V/NDGAOVOsCu1rAHuE4fNz2HYP7R1CowNDNaYV8hEwKp
dDk/Su6dTTiq6l20Q63LJBKdur1QFmJUjdfaZYQ5osJGtZAM7ZFd9LiRQU30pRE/
RA4IGVefWK6/jrtyjycUBE7BJULAnHI9oj9rZxAK/V3YNR8hDIKkytvGJBP2iKNF
d/IvYMKf2fI3+eX95lN2qWdHuHf6J4Rd5uVCOmWZsxz8KkTlszq/YOqaWhpovXHF
b1Fhbem70ZN3W6PJpnogxmUhqiNQHJB6bPduUgeqD1MraEUnUT4w0NSpWUVUuGh3
CE+NhtErNIZ6VNGotIBJdekfrG33IVSjoGDlywndMKGxpv8sLsRiDHvEDvP2ppkv
Ii9XD0bCa7vicdgog37VlfGtH7TdDiyZSXM8mrIbxtaexm9YDfFtuUpGwH7Pxk6c
62MN28PkpZeMwkFzhC4ejHT2R3OOBezMo5z+pImFNohKOmYBBxt4k2oynr9d4C2w
4+JJD8QPYttQgkq2wQb8YG95v8oN0HgPV0XAkbV8ZAnkynFSssjPLZObI5b9wKdz
KJgxOW8Gioo0H7DGLYlx+j6Zdlt8gHHzCvjqvMSEKfLRh27SR6xoTklglx20oxoU
YBN5m1c1Ac1KJG5BxO+xdUiUBMCfpaHfmnXh8YBPGf7Qs7+dSysjeslJciiwFG/c
Z1tvRGZRa6pjifgzNV8jMWtUhxxO4jXGJkOz/8f5+45y94H2m8yPBD0X49JUVXKf
oJ9aOETCFWdCV/CLFVnC6nrKdSYk4BMif7Bs36f63M3VQ+Cf+kpRnr+/PGLY21ba
+ZRqUPF2plkQZUQ2Riuledd2VWMZUMsXnOIm8t8pTYBbjlSimOftKh7dCbWAIZfJ
MY6lnTDCDlY0RE9Lnh73xmcfdOyUsjkwBo+RQd1uu1LoIbH1smCIBIxZbm5kiZfU
LktMe1x21aYLzWKNGDCcoyAFaf4KOsmD651ozecM6w6771VlWLKtdxFV+HU0uh4X
ytvBgNphnwU5jJJmVwt85MhC03rags8m4RSdJn2zRav1WwTwxqqeMULPwh98r7MN
oIQzTsmHKfd2EOAZQamYoQ80Aosj1141BWksdnbze2RLBCk4bwpQ9VSB6x/JrsCh
b6VsCT2wB+O5mB4QcbuxpFAuyBs3zFjs09Nce35xdIrgnk63dr/nF1joxvQv9TSi
Wgq7yMmoulHeKdSn4Ve8qWex7dz4iljdv5WjdSjWafQtXpUIFqwoVcbtmX7ASPtH
r3w/EJBQgQoP7v6k5zow1uO6o0QUKZijwFLbk5j0WXHUh2DMT5uGgG9A15UZXFbM
LueajUgIJ44m72DTYXrlFHNCyMTES8kc+BlHQnRLLHMmSLnM22UxUwDYm6hRJXq7
eD+Kuou0jmBa8naSd3PKyoDZ3P8g9jctZvIzbMfFfMwYvTPKccYo5NZHAw3Qk8WX
YjGpTEPdPARUnedhHFgwYD45qAlwZOQwcGFTu6kOW31UTb4cGc6CfbI++wp4g6vL
anPMmUmmHzOnRra4gR5OY6pmNBpTuAELBGg8EFZjXQp9o0YaDmSx5+BjmzndExcS
0T8b1UzV0mPwg4d06UBeV/uwamQ7Xj8YdD/Birl4QExZc3He4ZnqMpzNVMDfSR8H
O8qmaQqnh4KB0qDD9Yg6MVLmbdiwjsDSIQQAeeAHyUXdTPGTfwu5aWks5qIVrSW/
3XoG0Vfnz+eb+YmA3qZ+0QkQvwxfn/VC4AnjvMxwsv02fKUjlkkhN9hrt+jU/5c0
7FWIQB/0BZ+gp8efIiqeEys3ga4qjtt/SzeRwenNUCEPt2LTQaouKTZLFvk9dUGR
wFT9UBZ8IDkKVIdb+3t6mNH7ci5NfY1Rl3evD0EfnW6Df4CHW0SJ9/TH2Vil4gdT
hoREfI2JV0217dSnLXpKQ2uILFbaI4PHFRhoE+eZyIunM9kuG7K7Q25d1COt1AB3
XMZUU1lj/3DhCTBiiIyi/WD/Wmd9yL8uYxbbx12SI3IbpcfAC+udJh29Ssh/aLLU
ovfESdgx+yw9DZsoHu9vOoNi4yR0313MupR13S95l5+AYKuXs2Z3308D2x0ktuon
T9sB533LuczHCdY4+24zBUUY63k3cKJA5k4Gu9zCPtrV8cXZPdtq/dZ9nrvEk8S0
Ie5rci7TubI5esasVLQ5gp+sWz8EO5o+2mz8PFJ5b6pzFcMhWWo+VkqOgEOqEPu8
IoSXbjpzosq0hg6oOs7lUCc34Z9xmohf7SpkAT+0rNRZJ/KhazfMmhFoNWDRiUGO
WvSs1FYzDEorSTmQPxlmzpvXCe6pDxvFmyvmxzcLwYwUxnCjwWdOisvMkcHLE9Ho
v8OmkU75pdY1MFS6pvdMje+7t359ucC1a+fSZtG7bj4cI4Q6SvJJ20D7w2uJTXo4
qD1BrWWiz8Yzo6rMwqvjyvWD5qlDksZl6lg/7mnXsGYl8+xhOV7WpzgV/0HDSRaQ
sKrTMdHjpRvLRaFJgnHVVRF5c+SABmht2zAkvCXZzJzvLlvu8937NOwpIXSAkxOJ
BLt6AqdrVfis/py/QQA0zWIxsL6SJLW/jj/ALZw3itj45VD9J1v6Csvlcg0lEpcX
Cl2N+FGoCkl0nZ2aFheLQb8m+DnXMMriRrh/xfyZhZMSekpa9T++l8IMnx0671aj
aGTD0yR9fy/8HACdP6jnvkuk1S7whnYBteDpaooPZ7rRVjpTdNgsaB5AfXkhy+Wk
36SiZdxqdYEBVeZvk5zK5lOZ53x9uFAJ77EJxk4RzeCAC47ah4ccfNlvWlfL4wRa
VPwB8pPMyJ+8vAyKzVik9tBP4vm8qUWa3eAUGXDa1VGP9M6KOtW+bVWKrMv9rbkK
InBRm0NTWHU2eEJYQYB/4qOCnDVEFyWocXi7gT90MMOCb/E5jHMCzR0hoGdTPJwH
nGEkW9mhCM4S44PtYdO+0BxIB/YOuVMnOUs6Uj8liN9Cl7PxCiyuifUjIacP8t3l
V1uTFUL67IRTpiiwlWp4s01fzw/CY7KICH1FIHVHd9MCNAkg1msCRvXiaDsX+sOI
MQko5ZjoSVThV4GQCILVUC9p5qKCfY/RpJl5RG6yn14NefqRwexJUYMhrVzxnDVj
TSVu+ri0KUIK1zErjdwXVHpj37McWobxHuVl6D/2EMBLozKLOSziHsutNklnPFGQ
LvzeLH9+N/t3phGQXBsdChm2KIAz2QjbValtoKXTFLIU7QFvJ2yiozEWw9To8ewC
IJu+rKEy6hkG/bQSw+jUC+5O/IMSkDCKpMf2dFPG26SYwhfgiJsUpYOtzxqEQMjo
6NSQQ2CWw1cyQwrQHbXoKE9+HD0bJvwJ1WnZpP21IkGxfh1k5xn2tj2ZHcWEoaeJ
byr9FTAlybaYxuKW09hnS0aMVTdY+ZNsC7WclD6Ujz4V0J6LKyrTvWD0mRb+oYhF
4evoSLAg7QfrkC4UCHBu8vNFyl9WGQI8+7c93I9fCPd02KHWIDy4bZxr0Jgbp2m7
XwUjNhEY/+zFeyjMKr2BGMx00gYFeEUIB6B7E4pwT73Mo4+Vt8ysaKIl1Nvk6nDZ
mK8CsSsgVRBtK7LUJNy/CiSPWWS32jFsAfGD53FfiYoFHF3/yt9kWU1bwtLvghWl
YAycQvwO42PgzgA505m375ZBXZhneW51GCezGBQehd9U+87sXMvuLwZyrL9JaDSp
Ng16jLoOurq9N1wuSKOEfB6uqalNWxtLQs/6n8/cDSsUXqK7Xb0d03wmb7UMh0An
zgynZpS/4239qCpbpXyNoGpn+KOqJYmvnQrk9Y8yslAr9W/UgFk7qwz0L5G5mpfQ
oCArprDMfsEFVS3MJqGQHUX8f3+t+X0TYOdTQgGuyplFbPnqpWOUWtK+/zr9nIZ8
/0RaTl0F1YmTGWVJqSXvOh1MMYpZ1VxORv4Q6+0s0ClyhNazCs21+owHh8XowjxE
wkApR9HyYEvkEvvDx3FbnjyKDqfviIu4r/0HrromvR6nsxlmY0gjerHWgg09zf2M
31PpcN5AaftPyi02Mlfkdr/hB4bsKRkSuM/ZBynw3BJe+6AApZozV3jluiCE6nwo
8UY1fLsM+ECN3g8E6bNEGekp43wXuRFIs6A6APxvT4B3BoGmksnpyT5AID+mzTCR
Aa+4K7OPZM8bUFMg9MgsUUQf+N4vunRbwLQGFyo9OH9fYqntrYfLFS8qp4mJKdCW
aIqps/pV6cGB+jBqkYyvttSIo8Hd40G6Sf8znLGfCjRS4ojcuDG57y/2e1o1URrQ
KX0icHpM3EQhtBrM0sCbqPnhJpiiArMoNOGOMOeQG2f72GdimDYJ56pNjH5v0Y5y
YFMtO2aLL+Zb9+k66Ptw0qG7nL9ZQ1YV51buS4xKOUaZwPLkcBSHVSWqvKLUv/Fa
yCHoQ0mT3R3NeIMnLidQkKhnjmXWTJgMLe9KmCukTrmxSDXtynBR7Bb1UDxDWEJ2
4ji+LYzsL8W9EwICpFaXg2ItRZlYcNvuFUZo30fWEbOHzisIve0fxz2I72zs9RKK
0+M6JydDJA7GXvhEKcTH428MvOhtss3TkxVPqZoFIIhW7KJW3MoSsHkglPEGhYl0
sAlLEGJKaNabv+CiB4PBnxU+p5ORzL6OY4pxEEsIX+EpjDTwmKY3U85QdhVfTXPe
Jh27+tIcNw9oTxKLz0062HFbkkepzZx2wlk/uFh3DLcSYU+RDfYt82CW+ANr42Dv
l3ae93beHMRmsdWKBk+dT9EfoM+rKYTuVlTS4DttWsCqgbMysgMEafINaX9hyg7g
bI3+EM437lNRroERTMDLl0Z1KFTht3iDPHZEO30sPOnCo8z8xLF7i8HEdsg4MtF7
hWzVl+FOjyroRmkAxfpU58bVxuZhi5eQWpXSrPP7XmFq6G0103N4Syd1mKPz0yTL
rzmkf90gMjmQvrMqgJdKCf08YpPctBMzl4TzHzJxXveA3NDVuIMoz38xaFxP0l0Y
tzqLSDhAo3WqCxtChsxH4wii75BlbceYA5/4c+s+WDei1imtSUCDMuTcsFqysJp2
Xh42hk3MMw1bB/wzRpLTgT2hUiWcjvahiFMi3d/m0ZhMXEUpao6UAksy0HnhJUFZ
RN+iQYeGG5ZA2OoWH0mgWFM8+ClOP3OPsaEyxIKWyey5G3CGgfJMWidQBQJdZxpW
rwfIkzZ8Y3/ob18+Z6yfcUjAmkPUZqAq+AYE4ZJwHRMBexWV4Exb+NcKHYYpWtIG
VZ5y4fnsqlxUs5RzE77qtZcvOjdRRpBPMGjassbBasjiVvjb/tDLKQU4IR1GBl1Y
iK1Vj5GkrFt37169xuuHHZyWAfsEmFZn8oZSN6GuQDYER1gIPV7eSZSR1ymysWk4
40tqbR3ZjtidhVEqEU/31dVuHCMijO0/eNC1Rb3OeXvxdnC67H7HEh6plGxCj2z1
Q5WSqQmnFWYqkcr2553ctoDNdmjQqWrC0w3B/Qyr2pBKW1sS/0BnPn9UfQG2xfBF
JVV+s0xfcdLsgn5exgeQPFJmY8DUs0AWFIINFxmlbJ52EzZ4yr+UIIw+R4YEipIJ
4p39ibIEWtYq3aGgOk9CRVfzcV5QdyKUYLib4EOWBesOSy/tSIzEc4iXqVLfE+tj
drqIV0PJ86MrPid/9zSB5Oj6FTV+OX+8Mk75fCiBHtj7srBQyDrlwWnX77nHHzVV
/5sUfPb9XT5xOb8RVURTWvMHOBTAvbHz6DPq+CFXQiuUl+PQT0rEdUVdwxtQx5Ov
7IBHwJXw2emSY1HmNxxddqFUdVBo6R8BamWPW1V436xkvC5ojVvSoussWxns1yiL
vvZ/jUjFcCuLLMAb0sRP3QwNHigvaF+6XCaouZaLHcIlhZcMlz2Nv1FWt17c2HI0
/fHlzKuVtfOdDGVLiIwGUVLh8ZXABADWWV4K6jNHfLtWK+MxBCqnn8rZnUGPgeLn
/61413kw3oKkiqGx2uRi9WSKPPWeis+iNwiIngX20S/zoq68BKv79Lp9QM6TXBcn
NPUV20EQy6oLRON5he4NcMsPRKwddHBBvHSxn2FowAOjKQlf4ATu3WVfEio5UAX9
hEdui9LLvJg3NZK9rMEuD2SIM0S03U7epNNggLmMF3DbFH1Be44jsVmHI2AGS9MK
4yzhoUgO3CKiQQhY641DbYbnwLz+QlRewny/UBEuOkSklJppSGNXhB0tEFmskSIW
rPPayz7gIq/DU3XXSQ1QlYGRiYed9qnGPW9pPaPQ8VDdWNxutLKTPtmVc7mixW8c
Qsslu7Rq2rbIMK84TSmC/slm4N9oqhTJpYxUq4rCrqCGMkRpHQqTXhTcI7BE27lX
iqej02SmAF4QEV2a/srtJquuVfyKrAhxzaZf64bPX3TvycVdPSLYuLq2kJvH/s7a
t0dFA7Kv+KQlsi/um1yRmQ3O3HArP+STodkifvQISMmTJiAYA0zi5ldqJKkUCUOq
fm4vwbQSiMpyYp/K08ZZkR+1pFuHAFFMomoErdKkYjlY0v7C53Y9Q/Gq5a55PNCY
NCfS+K9hbD99p0x5zLmCDG9WQhWQbCoIKoNdytge5hZCbf3kmWu7adYpyWt4lLCI
NcBy5lFusTiT8QNBxnbjEceWjKKs7omS0vXPfaczYhxeDvRJFYSM7+S5Mo6cjpUh
B/h8lvWN7gaE/6aJdiqjv3pbB9w7jRcHsd9Kvx46QKKmb23jft8p+CU1++6+eIek
VRBDMvDaysVXZZZerw+Wql9//63DKZmTnFCOnsjBHZ3oOs30s/1pPGwv1cPQ3UaO
NHFO5OAb3PGxwSGFpzfEtMqEgLdAHtZ1OTcxYtOAQurpBcSY/ZzdJAUC3zAR4i4c
Wa5TUXU68h/N8+dNssEn50VcGvcGwPfOMu9BbRLEdCls2wZ1EqwrEx0d5ril5Q4w
qFtrUdiP9hK7MXOGp8WSqMG3CToB9cIiUdd7kxtWYSSM1Bo6BL7yIm4Bs2NzVTkU
9fo1UAYq38nj97m5vu06EUaQZIWRF/H0bntg1vR33bitYtodYU4SrjJie1GSVDHZ
kHV2o0VzeK4SL1U+mJOGgqPW0OS7uMh8g3cdt9VNy/s2u8wiilMQIidCmkdkXthk
cKI9PtQXyHfLFS6PEZW6llLYTiYe0IHap5OmncDbQCOp3OBiq9Lio4XigM8y3Tga
XK1x7u1A4hFiE4B92B+CPovg+G8XxZwWCnmu9NAZEDwIDISO2Db/RfJ1UGPSvUF9
co0Pqw7OM7YEG4rpssa2vPHUgbfNwIcmKcX1EF8zip/8AIs6zHvCIKM1EPIIFm4k
oX+hRcRV+X+p8EuGuWK7tXPszPesNEIXvlzHBmwiLMBEkKnxkvXgMPbO9FJ6sSz6
ufS4G55t4yqDGrwGpGG8Io6bt+BGvQP9hN03xEfJyoY+OY9wY18FkJXfiDJHFk8k
u1RwDaVT4Rt85oEmYJQfLZtigmCERz21KnaH/8DURxj3+ypslVIWFWo8vm9LHoLX
hrSKVf1T8lnpm4FZPHX/DNLKSN6GcWEdjIUas7Or4XXGvNfCZbBaqKzfAlzJgPLb
PuSOUk4AO9VhFuvqaUwHlzIjM0rvj8Epn7OSRmQf4gKNtq8fH0NtsgLORzxD4DmA
Bm/CIqbZoO+1hwZKOrgOEk7V6d3G3IgCKzsLdTnzY3SfTmK+9lwp+Q72qtTJA4pH
XcDrfXUs20uBGPW9zRPDgCg/VZ7StJlPw8nA6dbGnI6xcR+8ochOoY8g4xt3awf6
6Br4z/9bYcS+U3skRw3LFDj+SMhozV/4GtO9dCJ5hlUCiJHEQpCp0DXi2zBuRG9B
oF22sP6E8psbz2gpV4eV8BjvD7DBjow2ltvBrFRq66OX6iRmSeHB70d325z9Ss7Q
pE8I5i88FVf9WT9PrSF/kvEQXf03k3PjIJVHj7S4zyw5f+/svnzvYi58J8NUy5xR
8BdyYDEbrAAyQRaCjOScFyjgl/esd6nPQh/lmCQ2neRRZIqplQ7XtIse+jELHACY
F79NoH/5mMLZB/O3Xpwg1VJR/ZGE8THygBTtd8AJz7iunQdrJgmCSqLqPHhJXdyO
uL+A2/14FpMFcuwvKdv4WT3jW4KAieySk6LlwStgaMYtDUIQtnuauWDE9PbYKWJz
caOTKJ/S2+OkQjjl03R7eA+s5fhbhIdAhxKJSCJvOkO+C4ECGL9LnYLGyO3jSEaR
/T6tS059y7XxtiYCZCeqUwwmLkRAG0Ik4POnTNlUfn5sFYJ0PBqA/mJ1JbeogYpN
tDmxy7dW4AERDqQTUJ6v/Kc/wa7hJWqj/oOM4f9PCCIv1ILexASl7LPyObTRZPTI
Sc2nnHYseSje8iz2vxJ5EvOgFSL+5Rc3GhqXDXCcG9VhRPuCIFcZX6olNfMU+CWH
ygXJ7R8/y4y0BFF/OqbX2d56b/YWxWMQFJZgVZ74T3RwdEVhEANzvrxao2wAcqmH
YmtCbZ2ksaJv3VD04TuTxqJu4Q3G/vs5JtmNXxOx+mL/LYuVft2GkATvoYEAa7B4
fZz7KlQtWvEZo0p2xk/NJ8UwqIAsu8kfqPFQ+GX0xk4mOkTbih2qVVtOw331sI8c
UB1uZ/+QRZdXBbMZk6asKCCP4U02ACIANiwBXTOtWfMu23iXet5nSagEf47J107A
B9PLyVFm8dtOkG1ihIAdvtBiz+Lmh00EWYsJhTyohGITN+Z7CjdDpneOS2BSQ9p3
I95jufIXgN9UnBzAzGvbpuFXwVen5Iq6Xz9inLv8RmGVsV5yHvs3DlcSQGUDRsLp
gs1GolhkvjDmexIwV+wo24b/yFMmFFdTUU/RMLyk3dNrc8TT7IC72aUe4yljldoX
YX303P25/szvVXbCbceJrD8xRZ1Ypnb318uNuAtto4kGD+74mFFeQdqQtT3rObIh
knDRr9+l5Rv5OsFP7VOW/ApRNKqnRvaG+m7SKH3Xha/dZe5/O4pmK05Gdhn5JU2i
e9mmqNLfWw1yevLjs/MRUIrjvZYFxU9BgPTJ24g6OsJjyA0q4Z1+hqnTgQQeLdE+
7WLsJri9IF9kzkyRbaGTck32PeYlzaGZnrcFavjCKt+QmGcA6bv1BjwGgoEe7f2M
WrvafHtqciVez7JX+2H/70RpplGvM5juSxmki73Uk28jYojMKKy/vH2T6gA4umFF
wlt3SDF9qHlH+VAGUxiJHU7rP5xKOYuuj+Q2sTiTf4hf+cf2r4T5ZHh8atb23g0W
5iZbbdFhyrp9wtniRxe7jv0FfOes51Xy995gxeIHmDfSERDWajVp4EdZzPqPmUp8
PDZoFWqItuj+6gbXleEIsaHhJMYedsPrC+LXhi6aADvtUtBDnWBgppyETDsMrY6x
6+hZkGbL9GkwN11jlPoXW1vZ1iWCZMFJtZXV9GecBIMXaJq6jW67tHXB5orKrRPc
8BIO1nqJdzsYunOhpSlJ6JOoQus+bditXWBhMaxwwNDabRBOijSgCvS+I4hG2+Ek
2jp9ZYvFTyOuCPj9AqxH+PDZpgg9pefOHySZb7xCnLYIOtP6w2dMhCst+GlFmwRM
0pcPthmRNky9u7lUWJX0r3hKKBNueLJVXzcWhnkTKqLbwVpk6/rtBTj8I1KdCNoi
Pf9B/RWkLo6ywctmuzlzeE/STw2XVTchJOBdljlEnQRs9XRkNJcJoP5ybn6YIMxE
LbNT2kcWxnrVo8/2Metv7+0FBu6bQkCy5ZVtbqKFdFKqXIySdO4p3ndlJM1daR8z
ixrk8lC2mu/gGfKhIL+YnLgJslaa1yiNVSojUtsIUIcHzfj8AVzrc+GQB0SaUWg9
CHCXstPbliIZeOp7oJO1o4QRUxt1clZkTBcBgPLbzaN9wXCY3cO/MYMwsl5R0qjp
wIebo4xBu4xek6B2v6YlB1P3zF9LEeUKHPnZL9cmMVMj2rGJ67muYVukV3tWG9mS
btW3phQ8R9UcQvNJotbunarAwdFeLfEqtSmJBJxV/lpB7hQSthmbpvN2QvlPWB8c
yqPFZ28Hmbu4oZKaBLlLFqIcnUtjbtMMbc5CE5IjPuVCqIVgMjik1xzkDWQCBpV+
7FJY1Qhir4EG1JLQPqysz5QBOTU7fI9oNU1wpk+ID1f4j5YSLMmffRZvKrctyari
e6G6903a+PtpjNGy06pdvcGQ2j9bu8kZaLSlQ8IieYq2ja1mbSyED/xe/oqYMjYO
9Cpthtxx9uxkeX+5iprVOxzca0NuuM8dFrWIrDOo/+QWFc0NFCecP1fjR14JA6e/
OFWoNZRQDsf1ERYV/CEJyUgdbYt0Rb9JuajX+sTKmK1SdECWhvjMUcSuflAqNSwR
Qt/kHROxATkIGVyZnBmgI2UDqMlSCqlbBnHYKzOCmhwIpPv2/gAtNtU8ItjYYWQq
zdVkKu1M875N0/h+khsUO0ZbjBKUlEQpIj28JxlucjaLGuPoqhlIUT6BiEEFFn7i
ETJqFMra9LSmFPeOaYAoRL3OfAGJYkgeUlUC5mIrAxgK0IXtTULjwR3OYuW2YUeR
pKyWq8ExjZOZRnlRIdYp9WiU5JeMedTzaUY0gq+hYfcplbFDCFgfI0+3zNsl1X6E
UZeY9WOXKXNIR3spVgd7DtWLPWN8n0jfEFpjOf3cszqqvwMbVBMUdgzqo/ie0EVp
f+nios2QN30L0m/0Og17aDyordh5GdRptEa7cODGo4nT535XG7d9azbFJP7LPLG0
KnkkuQHbSk6kSHhKkImEzARVRWwcV1HJJYLrzkIMjA4AYxrKy9fX0tcqadOUIeEv
z2lRwF4V04VxuwfVEWwZjzDo9b2TBiRjZoput7YQ2VITJ4y2DRcFDdwXbijsUvXP
rDBn9VnRtlhmS4ai7PL61ZEJ+zjbN8raQVB2PeJGKYFjLt8QdPdrC5djhy04rPVU
54DajjmKBSKPY/wU431OLvgv4lGjL/5ljzQBrsye1uCYXqDYaITbjxn4xYVzdg8n
rhq2eTAMYMInaZWFveJzLqvNVHsujS6XWQ2NuGzRwKzrVoNWIORcY7fO7cby/Tr7
eIxj2GzvLmlFhf6UsKu3Eg+tgt4LH85imswBMTKZGMdNqx5bFCxT+GOMCgb7GqVh
IXoU0BExTJUKj4d46nNUAXeu3iRcj3Y7eGocXrmSZAY79E4mAWvPGbVt5tXVi77C
5UP/8Sfh/qz44Zb62n0fAvQ3GaGXXEHnzEZbw29lrsGAWVp3ubHOWG4Dz/mZKsQv
WAEs/ReIUW58S9y8Izzt6C0osyJzx0Q7NHAG6XITYNGV5ikpKKI8PtCk8QBV8lfV
+/y6frE7yn0Wt6iCP1QdvTmSGsumK2VrTV3Ug0eFOX09zhe9Z3D9LoqN9LI6JwjO
7KZtgWqHlETR7geHSC2TKEG33jd9ELoulJunLxnfFgD+cvBa2gMxxmjtGXol9TiR
7xPavpZy5pnH3HjU30xXxu/hmnpiMVW9T+qP5QYKMF4si9TEHf1mbBOjNC3cXBUK
Okl65JrgCSdJ7RN7B6W52Q==
`pragma protect end_protected

`endif // `ifndef _VF_AXI_MON_HNDLR_SV_


