//----------------------------------------------------------------------
/**
 * @file vpr_file_io.sv
 * @brief Defines File I/O class.
 */
/*
 * Copyright (C) 2009-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VPR_FILE_IO_SV_
`define _VPR_FILE_IO_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
XKdnLzNlSNAN07RGfTsValgLQAIgdF3yuu7YVzaFs1w6ydAZOLp53bW+mn0Pa3JV
uGL46bFDwu+o/J5DeMLV2bJWihZq9amGbKSvqcM4GkhI5xPxkecKRFZSshfYxbna
czB9K21VOc01tCzoRMjggVQEc3K3K/cMWidpm+oqBJkGFH/HIhUicQYqfkU8yWSg
J03A716yHdRaYdJxDUAoa0rhYoWVUTclfJ9eOVQbEYVI9RX4zi2LYpHDXULqKoEr
AtvBXggToz7UqeFk8urKQsesB4nVoIjTLW/5iz6mRH1JtbKl6gGGNn87nJKqkR+M
ssAoyP07rpOSZZufI5b0DA==
`pragma protect data_block
hu/zJU8c4oukGV/a/HZWbMoO1sITKnVU8Ch8Q2o77AtpQbTIwYIizx7UXPCRzIz+
OdWehN0GIeCWRokiwkAtIwHU1sUE2f9QmOtfV0w93Kfx71ipHbRkQd86BHSByHB/
M1qIR+d3bSkhjj3vY8WXPI+P9xXkt3KWFVFshlOEEIvzU2ePh6l+FJo1bDy6cb1q
baDCQljDLIf1THH4xYSdgf4vXg+boEf8cyuvAAR2EihBuPRt/QVjwiSGNNZHNBhg
NUySNR6WkXH+ev3gOmzMzQb/vYC86dYDc2jzQ4fkpPxAjCzv3APORJs25MJxf8Pm
h+Jqxs87UYzo2j6lkJpbn6CY3F6xPjqP8224h1QdhAsweSPZcdzfCvwUeKKbI4NH
sy/sw3j8upD0ygWZdDWXCg5GmIMuhYtA3dIuJk8b6eOcoU3/6tEWJDx7oWjI8Bbz
svL11OZhW8Iv5vOZAWEigq+nemFI6/eYJbxJhwMCULic4WzyjVMGWz+wNH8+IJ9n
vj9F3PMWEFNo71YErUnPH9VY8JBY97f8y/xNsgNMpmk/I+eXC19AzrW/yF75TODa
wrR/0UAHBG3RCvKAq0p8awZbTN6nQK74d5tmisQbnRYm2K0+f22XbT3CyMfVUsxf
EfI7As4K2TKw4E96qQCIhxjbMKJaDyGIAsRosYFiJnmSYzwcy0YDTJw+UwkOS+GJ
Yv6dqUXKeW2UxqdGUScPicBXJyeSlOsF0DvcvmmH0l9pJTlzTkzYjfSQr10DOx6Y
X++9Lzpto7DBDmhMh6SxPjlzUOD5LblHRkvL38PYP4IIF3YDZll+jXyhXfRZflFj
NfFCApJpA6rQVDYgegWASncweR6nSYT8zlK7xiRM8Q9Wo90PHQgYNqSzOxUDtHGb
/5r7A86kUZ8SmI1rganJbzs+COxXkriaRIB870KduATGj5O5oXHXk9hdMNLZvHKX
E75zx1T7cW3sxOoBjtzbcDpqjfSg4gwXhQntvJMbwr7/NeR+xGc0ThmUCYMzWOND
2rA6BBoTQh5MSHGPeFAEXDHmWl6bfTxhxUWqS13iMTOQLFBlTGSTjkM3PhFtFVdx
CkE7tpZenRD3IX+RiVr70pOjJJCyCy0hcVeRThKYwK3LixM/GPEwt4E5702va9R2
37fDF57g48VI4ZaqV1JSUHmW1WR4+0fUvVdetvPAHt6YoYde27WDkdmoJ03FMDyu
ys1d8W5Vdd4LXTaFJlg5qmO2vvQfiXT/LxtENiXDkKmL30k8e0PXRy1Pv338V30F
UpcWvsR01AS+GJsJp/rr2kpCfGCm6xOHmEBjgdMMM6OnRlBG4Z4zhMaka8BSrK+b
h0MLY1g6qpsaAmaWPOevPu3cEZm43UzXOp8zrwUt2p5JAiSfkEF/YL/GV4pHjxIi
1qDRsQl2IVONHXsnWYebLUgewuVBkWdQ+L1sISj2qJ0lSEMn/TsitDsLmk8FKRv9
Dh5ACLa88nqUQ+QdbQWqSdr2JapUal9pMEj2/WiuaLk+rk7ajkv9DqxC6v1hCS+k
WJWDyRRkEPSswyKQx9A8SxH9mYLM9w3xBTh+av3YLKJImnFD2DcLh77BfImYLDv0
ofNkvUTGaSPcKPYkphScpzGGucSpa04FU5g/eFLiB/L43bs0abKqr0oXxv1ySLl6
do8B6JArMmSQE7N/GZ2pFNjmG2xhj3JPzssgnJj91jMSCqYktsVFEl6ifTIfUmv9
3pcHF9KsbHClrMiDZ938+VhesT1G77BCdDRDBU/qRZVSBUY09bB+gb8hnlDG3WpS
/eDNPL1dJ/tksTN1oo/XXtubgx5taVtqJnZ7Bp5EoL820lqCLtgzTj+J0g9oDkSY
iwQTEV/zPy68ZJ76YiK8lc9h33V6Lz19Np4B+UQKayz+gVfBfhDxVS9P1ZMX0epa
80x8FEUR2vGFcscEebkcg/RBGuws0gvYCI7guvJmJDdfJnqSAvLylx2JWtCMVo5c
Pt7hgEHqeQWZKkBallRHYt309ZjJQMGPBjnSUGRZ8vSBOXgxhgOvN5Y/nrTo9nns
gaCxSOkBmJlCcK1i4gMzqkVRpSkKVaXUxMDeblTLWQAQL4oABQN6mt0kpL9yCK9F
oAPwenHowXVWrAbf8wkhbAG494JdgnMsPGTJ5Ca3vQvRaDjwBBUnDneSZioy6DwK
2gOeOAUcSSDffr+/LTgvu2WQRcA4qwgEoxx+iZko3ZgHwRxeVM03YQXOJmHG2oB0
reSV/TwuVvpjQFTQ6dea9RmfOHN1pKHFh4QxW7nfewVrW2nW2GxgnucPaUCuMtfY
A/qhdlInI9x2xiG+pI/yM7vrkI1SwyalVBIZ3f9J90kN7qk/jzgLpWVePhAzEhAl
/UTmanywkQOCMZKabMUDY4iHza+SP9tx0TNdNRm2eTDc7uDzGg35SIJG7nVgLWH2
NvKBqbUzqVHfbBZsbtOV7g60+QJQAGYxyGR4W23nMXXhsGKcQGgjffdsEHmSjpfM
X+JKDa63oZTkOpZ49O2Ley5lKMCwLudSSSVds+aqMYQgeYms/lSHB0NxSeVb/8ux
bRrCNGhwiw/ZmPh44tUH5/4MiaKOa7PuYAM0bCgB55MJrtv+6avk3u/5f7Q+lZvQ
8EmW7R0fVDOSS5fIIBuU2BVagAFd6HkRDmyFYDuiROSqwWObZ23kl4XB42hox4FJ
V80yygSekgraxLMjJOo4TU8k6NnkQpHXhesQFvaAI/fuMuRdfo7ybIinW49UAhjb
0+Vj5cTy623Ls+WX4Fv9AEHktzx9b/vskSMwfAFAvd4+a8kVhzs6zzAl/01C8AFK
OXTloeluSfFBKQnV7dap2L3vVXXGmqDK1F9aJKiJw337rH4zIPGrOX7ZukCvSXbB
NSIG4PFFSohA1hTuhLvA/CITfwE7F0M/6wnqu9yLV7jHnnDCuYFPX6PZ3JjAOr4B
XFBlreYmINd+e5PCFSEW/EykUT2s5SWKpVdYy6cbrdktC/YLfwfQWMt9Q7ilxaVi
dPRRvbDt3Xab1L9n2FbOBB/69aT3FOggUheJJLb537bdx62+xZyUv6K9S4M1FsvB
suacXSj4Y/P5SlTXgmfJAR5Ar9BJKn4GzAUuQ3jtyQsRGFpSo6G+UQDH8Hs/encl
mgL002Z5eZRh1a/Jt+ulXOiT6x8RDpoz1S/QVOZdiFFVuYSFlunFbM8jgByC3k0u
4oCyBzkJFwYDnXJhLvBR7m0EMmpGFvntW26/wAKxa+qrHePS3tjFsDx0i2n8GctB
H1FiJTRVzJjfQEdrg/uUhhizmt0aAyv5IcZeSlM/65j35FQ9EI7xjNICGPB2GmxX
95h1mbktD6v3Bh+TlxgajgtT9z0NQC8oeajfNDCnAHlRRgnscGz7A2Ov0aYObHSQ
nKL9TMsuWjW+SFWi2ZH3s3lmbNYkzP4Dfp/bQzgYSrO/lKGyxwHnZy/xyZtiFUYe
a4xdVQ8DMms6ysz/AJOMo6rEAl46b6A0wwSJXaOSxmAqe8YsJgAh85wu4lcTh3WB
3S7A88e7seJ/3CKNhNVhmdhpI8zB+jRJiqqE8cn1nHYzkwh+YZyUF2LFAt/KFLbg
I6t1dbo2YINKtb7Fync0nDfBvyhv23ZfqV5k52HwntjNY3v/wnfXcdExnSWUlsGE
tls2HS9G6WT4QC7TMt+ZCSGWqTzrr/DQlhC+ZRjD3/Gz2Nsni1234JhAmWsgdL+6
DXQ0EJr5bEXG553FGENFqrCKRo1vLl9Yqe1M4j2UzY4sIQboGtBGjJ7/cO2VrPr5
yBk2MwfuG+VW6jQBqiYkvIWnEy8gp8x0dfvz+7PSugsYN4zI8+bzJx3i4dGHzei2
cn9MiAdnZ7I0PPnWl83izlojK+HEcAWivTkc7AdEoTin0AnnO9JD9aW46rkif59D
hS354dDdU/aglYRQTuu2ILAkW/ukUeLRjMEbQ4/qYxJOuSlY389NN+dbGhrZONNk
IJRZjPPq2mqB/AOO68wNUb94lJiUPbHFOghxzvbV0M/SswDGDcndEfSZDahhC7mg
XUjNGpVJ/Ts6WWvgXOkmPk2RHJuhbTKFOjFUujjU1dUTg80D7+IseGBAMR5kjmrh
hiko4lUtzMLpo4bg0Kgj3iQDMUJI+fQtw3qgSbyDhXwjshX9nzQSNPmVh5GvVbHg
tQYL37TwKTHIHVMs45qjoHymAFGPJ1ofrpJscWDlUZHi9Pgh/6eNZ1Sva9IaxOBh
HB8heK2n8hQHDGRZBQPVfxpBWyUZW111MLk3rbrMWcRjtDZDBQlPY7FzIdbcnhr6
Vy6l5HWkqq+AV+ixoKDGyCW3PD86sTJRIfcj1acdf9PEj61wJglUCm75fnjny0zM
fNOO6cDKMH0nhpsi45WWZ2DVtJdfncObT8wcu6gviOLvatI7R5HlkKYR/hjHxBDr
NUGwS/edRvOIVs1cMb/T+hx85r6MC6QL3DG8sZfwTQVd5WI0Ze1imjjJEFYU2NPK
5kQmboM1SeZQVO8OjKKcZVOKKxrFeVWvhTSPU29Lz1dnYZF9QFG70UknzL33fVlw
I8J+QPGQY0Qku+FvMUh/5ZoTiWf5lif9DypWXhgVwehYcYAXW4l8N/0qWZgePaWz
WiAGq0F0KMbaNfaKt6dUA56IdN+fyqcOrHGZSomcEcgVUF8Bf+W/CpcadQ7Jpcl5
KmmFPIbLHVy/a568rwWRtaiqZY7g7SQfiZOcR8fb5qpxv9n/fSuHMIDUiUvOSunf
lsfQo0aFseS5gqoYQQfz4sAzwqYlAk8N6ewP+1IKQbPfa0c7zBjVWppzc5hVS7iJ
R9q66kb8Bg1HQolxsnjzLJ3kWo8nZoM3dOTI8gJt3zsat5ialNal2gzk+ws5w137
Hg2tnP89Z+kuHCEsgRBeB2x7GbaH15vnE2NUMtAuKq5JkhKYpR9gkehAGDN6hYH8
6/3BWmoCGuYe3aeEdmh8uWhXkYhFfRLPHM+KujZxwn/ZQm0S3jr+cgjQAvLs3+/R
AgnzFX0QQFCCrZ+UN5cTDOvIVr8xLFa73A2ODHvJ1zpLECgGit09QAfZAk+eakQ5
ajnVcmi1AlKfDnqLyv+00St6T1V6D3FyRZtbxhYQgJI7Sr7kNYHNmbVIBfsGy2rM
AW1dh+zkDpm5oq6e6HUYmLajIjSKglKR9N+Y9WOCBkpQMShoYW1oUUJsKLarL1QI
N9tRiXugejqiPd5LsQPpEdkoF/04pGKcQ+oZgq4qytzYyar1SDrm0jrX7Wj1bGeg
VDrZv+qBajssVqADxmL6AfBdFwTCKgtXNxd0Ga29lDr8gBtZ17EgcUoaCYXjDgQU
0n4bKWAyXP6Ta/Gh3/iAnlcJn2orEUQlqcZUmgAuHZaU4RG9iDw3hC4kk76ne5it
mZBO7oIwRJ+iq29X2bfEdkycuwCDA38SVDpdA5ZPqjVcRWKELhExYiHEG5mV5q/2
PPzt0BxAPUdkP0/rNhuFZq3OyHyzRDg8OApyRKNkbDlJmHSA3C242o2n5JyzQfSQ
kWgDhhOWwvc+P7l5mX0PtFfEPQ/38NwfhKq+0Yn/qBQtsfEkz8Q5X2UU5tPEY8oL
l2ej4JO4EBPblIOQF46p0KbrQAh4QNqeuus3AI0wERWNhKfECgCAAT4rsk97uJM3
XMEtoYS1R3EiS6yEHRF3d9+vekqN16jN4F3HWN6sFYsBnpEY7+RjO2Uy186d9SNN
43/2KngQipGEAQPnlbDg4uDopKT8qVLXkP+loiAYSgVUaD/mXagYSEToooJcdpTX
IDdLCJXXWGWgYpAbYqtHoMO4bm+epA9pjqYO0Y33kLtWZAwfLM1XLXv1ep4REOI2
zCVxGo8iNoUb6XZsRjIb8rG5rFSLd38Fm5q4l117mVxri2UkM44xA5hQvPLmyaBJ
2lDVdBbOK7Fc9PCTpXP1tpgkoao56bcPtB2Sr4rSDcMpi13C73XPOjInW++xvyLd
s/eQaXap1x5hNOHtuVfo60DwTpa33SshazYYD1Ihens7KnU2Ioe7w/2fGv5HM2lD
7jJms7S5MH4ktWcqPskqNaxVT4OrAh+N5L+JXByl5j3F7inDCYQmRnyjE4wJhc6N
57eNzDEORA8EYykyaF7uL0RKdUWeQdoqhEdOpFPjY7M9An5g4AQG8qGZjb0/5zOm
umaTA+P3AAqiWKLhVDSIhpLQfl42JPefcb2NUs1576l80d7ZFhYNAaWBdnk6OTAb
AU3yOJI6jAlio/uTzaUg2/iJXCbOzmlOk90YNRoLAwYjmnLjsUS0YLJs7RvbnYXr
Xk1lqyW84I5HvIiGCE4wOmCEGTf9EOew2NxjGH3mCAybZLuXnx4otrSXqtbDCW8N
0Kmtug1RCCyi8GSbu0r3Rlgeqb/oXIzsmQv9TkH+Rk50g5Na32/6VWcwWuj87C9+
1AijBqhLzVwtmsrpYQLH+WavY0YiIDHJekpq3Ms9eV7Tzll+MhzvmdxnDw9uM5d8
6tWocSxhNN6UCu/IHxxDp5davUbcZo3kx6hhLcMRBHxGzjis3FyxKICnrSl88DyQ
+xuQPd8lhxZML1zQNza296ThbhRA5npSQIJm89VvXx8=
`pragma protect end_protected

`endif // `ifndef _VPR_FILE_IO_SV_


