//----------------------------------------------------------------------
/**
 * @file vslib.sv
 * @brief Defines Verifore Starndard Library.
 */
/*
 * Copyright (C) 2007-2009 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSLIB_SV_
`define _VSLIB_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
VQB+7Wb7pP4NcMiudfVTFsBDBqF7zSS3acAWqjEkE1HaHWX7Nubcpgd7LwrDILf5
vwfhzq5aS3cElqosvKGLjjbFHjQy7MRychjcE3fGsGkwiIJk+nHvu8bmThIHi17J
OY8CioaEZCvCbCxxOZYKoJkpMzkDpkS8DGPI27kiBuUCqpjRMVf/swvEioDzc6oG
BNomQC7LnjK2RXE99jpFFxh226yIYow3jxxEzS+tm8YB5fVkTFp8neJ+JJR+YdAY
s+zRWr9ZQlrwpOFJCWkdDyzJFbqj3OAvzd8k10wfahyR+9kdnFSGxK9C9Ok0wYM8
7EJ3XoF/BO6b0KOWJu6xvg==
`pragma protect data_block
WfTo1/NcN91F8mOcSXqwkS+4Rj1P5CDboHFRIitAp+iv/CUtQ0qOgmwff9zBvBQs
en+/q2xL4mf2uSzFsCsq4Yiki8roKUDmRf5uCI6Dam2+7A/F5jvAvbMVms3bklJJ
biwlNLObrc83/8amwRuqpQ4Xo2iXpXi4UkrVtmCtzqIYydM216jZJVY9zLUUOZ6U
H25LCbu8W05e9bxKHaLk1ur9iRPB1/rArIeSA0LnXNT2uSiAy2aMhVbui2KQv8u0
S93XLXo0qbFy9iPtaKLfHErcP30I8RmVjQa1QYpRwmYVR3PRx1KtJ4t6+Q4g1JOg
nko/EHpVn77KoDUklfkPMisz4X2AsavLHkmjR3WOywN/xE0Vo1mQ/8CMWCLXkoy4
Zs3vLS6eJ8Hw87lx0xYfhgn6R7+Uo7K2nnl/5uiSA/kDK/Hw63OoonYgV85cyXAL
5me1RvWt5jYT/Mk8cVNstLJ7ChadkABtlyTmI6PQ6MvX7EncMphybuow1lg/Rxfv
/0puDvCjBwNiQ96qFPuquQ5RefjVti4BA2EsWIBbdciI1N+nkBqCYaxFDM+qQEHd
+SHxwYWZQAj7GYmnLaU+Pv7xXO+OSgepERbwcNd8CbX9x9RqcqA1hxkIwKJyBnUD
U1lRjgMAg3jV/a1mjL3/eJyqupNUiPuksi25RAcLCnCxGE07CFWvVnJGSmvwMrpx
kpyXnJ0Q/FAZNdL1BfBuaEZDhNZmELzVppjX7IJaniGS5bPiNeV3P6+ubrBwtZNa
+4LUwhPq81HBooq1ErZOeVrzX8p6EpcqTLihgJCXdlthIJ1xgtaB3EJxedNymZnz
D4HOEB8Fx4xtVJSqXXZHN0CiBZpgIKWxZftMLGQjvWkX2Zj1IjVGu71p8EOpIDda
V76LWk9Uzh3os9CFONUt915sKj3rpfGblzb6aYNGtRaRGL6ARrafskzFauy34x32
DmJ118SZx5TiKR86i8vfaBIzLIrRaKYalFSDOeQBYkgS5BEf8HrGA4qIsS+hgkw2
eVdMHK2UB5fReFUlTmXrehCAGqsNGq58z6LfET0qZHYfKoR0Udw1MMk8L9hEkoiA
M4KSv6RfOuolUwlggovBjkM61rq/L+ovtJvgRg4ITK7OHVz7If3EnJoWxspdvKeM
52kv7DLRF55imI/QlqWoggvacqXMBpgJuDWxGhEWILK8rsLTvd51PQV7SzJQrqnb
IgjAZMx9zErJQ1pedq978+uTInexphElw90W3uQNHU0RVRmHspVs8OJLDPfIvEzH
FVSM/9nLdRDgnt2v8X/979FFZHrhT7VSDnC6Yw3ksYZbAY5XwZ2FYCBN5ZcUM+Sy
rHVAHfG4i5GZB+ONWMwyOAj2CVCyf9KJSuA0fJjK29XtCTPuuU20QNFDXqpIgLtY
QksJJXN+DI/6DiMme6NyjPYG6a3IzTtJ9aN+pneZzZq4RevFmlw2KSXzBz3HmDB6
+/RFqd8y8OpizjIgg1+oPQOiINQ24qVIUWzaGWsPJtvKzD4eF6UhTYzSMj0f6Atv
JyrwIkxyBI2hWsB8XbPOy8L0hC2VgyweMJxeLcM0MnwIytYKlXRtHu7MdCbRJDD4
xN6nAuMdM6/JtRDXly0rGl4ubNDBO5sN2PoW8k7hgiSAuRuUFgrPR15l+tSyxDIi
slKc5ZEM0Elyzu/iWoj9PmgFu3C/hrQN4NO/BnoHsqkoVq0WsM69lsjhxH7Go9hA
2XA0YeBot15I25bixB99EKTvk8lLdJ7r9+QUgRG+POb1qf+lAp28J9bn0LMhNs5O
6NgKnk0PyW/ca5FrFoP730P9ogsOXQijQhP8JZRsl/jTqLgFaglFyON6Zr7dQD4P
kr/XCuy7qVu5YbekslpKepEyaa3WIpFkKrDBgNz5X8GA1GaBRqGll7fy7cvMgx1/
MwH+MmA8WpKPH4AEqfrPQvMwNqAtg+ysu9gpTb672niga1iYQTOzHoVKYDfHzCrr
ZZuYLegO+ThQLO31KiaPm8IwoDAkesj/wO70WX6ryM3m9iXfuGzZ3JQeCz19IXYQ
iXvEeIppukN3vtBZwgTcPPSintvVktBJN+5knYrSmn1cHyS5bcRhiJ8bNd46U1Tb
A7chluNXMlq06EXQ9ayIn6Np0DhYGNFPOp39yfbrAL1CCoZ4KzIEZS5zhBV685dr
gf86uKCBQF543qI/KEClf5YP1PoENvrTs8HQ/h3uPzOen8N3fA1bhhzkAC9DgQLw
hAIiQfzz2KwVRS3GWAC+ijqlbzllyGjz6ifb73Zd2W7cXalyxvoTKV/teuFhCZJR
bMPe9AOmfV32gzvcFTR+YVntt5pKjn8sfZtDPBs4zqNDQQDTTQUYl/yB6VEOhBwU
1taz+vIoSVgCpR5CKtKpf/nzJb9pXHtMnd7Zbb6LwzaMJ5RBXyKd9rRcEGp5Kaik
r0nr2gU8o6TC3d8NqHYTLTUktUUtlwIF7wgMSmvBT1BcLrHPgrHmehxMum8Dci75
4LWxJL5ePF2lJDIy9xJR+6QmgkzRsGSiuCryQnBmhlEn+8K0Ea/kwW0QM+0w4fov
hdvmawF4gd4xVICOBm29JLPWXuMJjkxCuPM/lV6K0bRZjh+B5OKQBCLoCpDRBAjG
t/4MuvD5pMY0276RxLsU/8ldO5IlprBZlgNl5KNKIT9bjH3X0pmadpfBJMn4+BF7
e4ogdeO8VKVg/ns6gdButVo8WV5+VuUdfe9d1inDroZVWLZ7+7uekuo42OGcHC8N
Nfcn7/T4WNrozzju25nMqTRcRflvRpU5Ucki3UuMN0Y3PUQEzylb2qZkIwnHBlpu
at5zyCoRCGThfcBbD7VLXur4l8QqLBiJN1xnvRkiwuzVPAW3g1/JH5OyH9nxlhI7
LZubryx1kyd66bNQxVqBJFgkV54oF1aKNBRQkGZRYS53rIP4AH+wIn9Q9l9CTjPd
coixTpSM+khNj5HiNZgrXJ1kbZnNB1L9i7q0icaGZ+kk01Wl1KiMbe7GrevoKl8K
vQM+pUSSGCq1mHUMF6bt2J/t29eNDpMb+Ycx67loYK6m5ZrlHcvlA2VCVgda0bc2
UF+oxOuUgaHQzC7I5MclSVngj6HcLScZLc6i0FuD9RzYuGj2AC7wUSY+5kH8A2tW
WizoxBqPSqYAqQehquToNObPCpgOBcAQ6vTnYGYdPfhAvYCfDrkcwRZEFMIUOW39
25sddMWh43j7NjCdtY7nyX7gk29H2XXIX/3MngVLwdKXSTmfjWZFgh0IpLlC/Ont
c42E0UYi0bqSsXrk8b+/nUh/GDiVSlbFbqFdcTZ2nc1C85aB2r9hzot1l+/nYsYx
+At4Lr8lMY/SoVnljH8DQan0zokyF46uhuIEw8+k0LdtLkSGGgPX+OiMjqkt+hKN
TWw7TnthrjZ7go6ZaqG5/njEpSdEK2qjzgiR1mhU4D5imvrJ1BCozRT8L0iSt7xd
fZ6brRWIzSV9ARQFs5DmRajMpKg79iTR1TFZpU7JfDhYZydYPpKTU4/akHzzXfjQ
XYJjpSq9GSUnumXLW5KRrOyfw1Q0JDqPvDmS0gW6gvnUp6nMFSqdC4VJmzM+vNYZ
UlGiM65wXmSDhNxdEXT6/SuaXaWE/cb0/OgnLLVnQP7RgNWAdGytyOV/ovcsqexk
pqEaVx2pRbNfebWOUCQlSCdLaSB0r5tta8F914Wyt2TknacgiARTTchWO9tphztY
HGHoclNan8dG46W6yuQCjHjdIAulBDxIZaHyKljPcI5UEnEKlVxP7UoV3i68blCN
TUa2iGkMUbFNdGLenaeRd6vbRsIt3rvztLlVh4xmvvR7BtyHRMmOHIh9aNtCYYAZ
p0X4cxes9Asdwd/xpSujPJTEYvwQQeXGvzww3H/5/vcrPFWbHUHIwMJFvynr8B0c
fJ1QlqKTpFet9IhMsjrVumw4e5xkLY5a4+uwmRjKjRU5nGF/7NDbNG6hKN+PtUDL
cykMrjx1DQCjUxM+8Gy8BmETi5KkeJqiLvL9SxfG++fYsY7kEHIuu+kKQaD+5kyc
T6bq3naQjIwCR6s56Yb36qlEUbj2Sj2ZMZcT4868xw157CCLhpUI5JKePlXWEkCY
h5g8EDnXynmNP4E327vBv+SKV/x8gCPRlPf/ad04RLXjtKdEIxeq0XqGTes3SWMp
Gs+F2oLE6GSSbFX4PdfM5cyTQ8d+eVGPduYyw45qMmomJ2AKrZa3UnW0NtgcNFS/
G+QtWVnmVzRfv1m3c/pj1/0fhk0XBWqmDHsueSpe4gb6LjHDO62mXb5P0IlvBSTu
/eZgGeA+eovayUvndqStPVFrs5c+34/hh1cTbBSUh3XIzsmEwrksT/2wsA2vJLy4
zbuU1icKFLiwB7DDtoFgCyvhrKwjgYD0i+jsBM6lqh1PmaHQV7M1FV4kx2/LW79G
dEzWtSAdoZF0qTMdtEib1kCcY0b8zFJHSjEcJ3koySwaSuYB/L2JaWsYpZfFqhEX
QW313AgVNx0p9AEgI5mDe+FdoQKBb71lO+ovoEvJN4iteYD0B67bhg1bhR3Q7K5O
oCb2YmjXgqhRZG1VrkgYsSLEs3KxZi4nZ9znfxbR43flScdcwcw5qc/2pKXtUba+
XjZ5JnMgy+eWLv5SBurUIq3DPbbMTvNkPxK9Yfe/4044vfBW/Zi0QUmaRsaNdoxf
921VNRBox2S/nkLnKa7Lz3kXz0PfjrHUVDgIKPI5vCnKmVAZ6f+r9RSFeIkbqFuX
8RPnhT/ZiQDAuUZHusvrktsgryAb86vbYYmSRaiXYJis8fOSYVczrCDqqaVn4x+9
OXd7YNAqTiHr+CdqtsJOvEZFYeef4SrYuGj5UiHl9qFfRGoYHehNr96jIxA0FVCr
LPqFQuOh8tBH+DBfxoGtEvzHjpvSJPjDPUnVns4Yuz1hv12h/PH4t8TL7UmISw3s
BRGslJWGr0Q1hiDPSue8HsHNDA6LwqKH0blyDrYsEMVIh62Rel28slMsP4EJRnob
XXqxVIRt+WfsO4J236EWsshKvJiT+cL6guw/mkVKkwav6eN9riDVTnrL1xJHMKPs
JvurYkWMzEw6o2cJH/FMkFuuoE1xPczAC1Alj+MvOsAh2ox7g8TmnAxN/5NaE+K3
g+R+6ANfat1V0OAl/fJufJcBqFZh+issU3AljU1UgGDJNdgqGm6rtZnYW2ckpHd8
NZzxCz2QqRXhR5D4Gt0BZfjYoPjKWMp/0QT1qrpBkwMp+RYcJU+uFjpX5q5yQNHy
wWW16rOd2GiSURbuyKAlBLvoBLLIMdk1Syq/rzhxBXF2HiBoRWpgUoWFCjPChFM4
flguadt7hLUukWcBHdXW91TQfueI46Afht0Oi6W/UDsicCaOKo8+cF5yGo/ajkLY
KHouhR6Bbd43UnpBSbHr0vRvFxFGX5Lv7LPQtukE2dVNMZvAERgrF19GCDX9JGOl
oCGVMvJASVFuJ97fz62a2jaAbKM6TQpe4SSc1HI+t2oHy7gQN0Z7KuI62E/lXuJw
Oc+J8p+3LBXbFAaBXcRsTpVwNWNmiI46zlQW2N77El1X+kABcZwR95iWnwJi4F3t
Eq+gLAPIeTWp0g3f90j6d1UKmnQ/3xPAYPFLlS7UDaj021c3FAhMAQ3/zx0ZZXss
ZhL5uq92zJ8M+fjti/Uq/DnbEQIFsiz+TmxOxqUOeWDtsAdqLXC1Dme+r5FJtKtU
SSNmHziPkTyF/IbwTnv4q+6932VOGXZ9sLU+GRZjSil9tB65Z2dFX3gHq42sdBF4
KBodfrsAjstIFKjDSjk+KILBl9+N70E1vVfqogZ6Lrq6pCN4OR/D95GdP8K4OCkK
ZxZFpWa7dxyBP9dRdvu6n0RhxE0yYvevxGmoTbG4aVT3vH3L3rEqOndsbBoUkhJ5
38PB3NL39M3uGBrpDs6mMvlWyrZAFbXwhLd/MQByxSEkcKw3YOo7X1UgKYbQy9wl
LSX+QtAij1a49dbvvgjF9Ol8489UBvF34PMbJHFjpx77TSBkc8SFkO2Qg5jz8kFi
uRBHt1ysthXEebK3HkcBaPEhPLCoCzhtsl+sbOxt2J4ccJdNNrnob0YFd38EX+Dm
i7nTZGcS29OV1EAnS+AjD84ovQG1ZKWHpWwQJGtJLvtgQNSdrtTnSOMp30xJSsEj
4xefE7vFs01kgaVL+k4+Pib+m/KeT/Fd02oC01PwGSH13npzQSFjEHEG13vTA+IE
To+swGh3CmatlYoEWsZQO/PuFs94M9uqwdhW0p6YQNlwU+46Wk7PEP59zgvAW/6r
ax/fFN4l09sss/nFjt76Y3UoSmqwegdU2HG0QOIUvSV3Hi4c4xa2/WFZNnps3hJ5
yI6mEXdjCk08ndET3e4D/LmjUJMY3iY9yj6McDeoBQFEyee0k/AvPjYo9J2m5ZQI
QD+WkTkSwDKRGPTVTYYNafq4VCKRfIL9E/VCuIxpP00oKvYo9qDDIhL37u2hGc8l
5lF97TZ7L/rClZUdJugRHBkDWO1i0Ii9IuJzppIBckVNRQFu/oDHKFAACFtgUNQ6
H7mmC0wi8O3hb06JvnnJK3J1RBLuORONWHjbX2MwopgzABissXjYAjRnsCTmpxk6
klvd8YN8r/3IXiVsohSKeUaN45FlZPsp9Wc5/nGojYOfqOxgiPXBslGdnIiT4iyI
Qss+7IebqlZVNGLAuk0CFBgrz5hOr9uMEWgVJM28suu6/+Rz3MOYALgM6NUqcR2k
H/eyKcQe7vFEBgRTMxNoKuKSbxbuBch/Z8oODygxq/wLgb2rGH4rgAA4i+FbKyHs
A7BQJ9RtRuzJHu3IwYydG72MH3GsA+dppBK+57mnrTQRNhq6HdiB5G5jLjSHOoDr
+vImHdvyvM0Ws6h1dMGCEe9Af6RYW0YnR5VUDUfvLX1GB+wR7zzLXtioexMk/hc2
Q3csyPb7lddxW/lCzVzcA8kcbZrp5Jg5LS+TNiGteO22dExxfo/p6UmL4yiZ+7+E
2skMveKFaXPDTBzp11M4qgtPR0q4K5RNWcLc1MXNpK6cT5NusOFEdsOi78aLyBKr
eUC4/Px+hAPgPPix4RkhgozLbmF3B1rKnH0dRhnMOrpgoqsq3e/46qbfcmeGUZ9z
B6cgy3pucdZLvmPu0tWieibzKdfiblKRTDR0YXq6rP3N584edqoJO833TY99ACkm
t2PetMjv5Y9jQ0lf/b6TBL1p0K4OygHRS5uEDP5wqDi5SkRJk5g8jGwf24TnDYKN
ONVMofyFX9i96IIzP/8XLlDQ/3J1LaPzFQXkltCyw3WpHL7xU/lwO5ifdEtLWBD7
xB3zODos6/H+Kxvaupvzr8zuK8Jt9Z0/fLFLJ9IxvAAe4cSLYuLb072Wn2rBtt8+
Iv2Qo4mk3Tyxwe+cJ4Q27wTcVdQsF0ZFHIdqvc2iI8kbLKjfhm0NKZZXE/HmwZ5L
6lJUoYc45f+C25Fp96bJKdI2/iVtK8e5tqsmNnoB5M6N6SyAsmi/Sp1XpCvn+wxy
+dBMJwOtgj/vExUKmr/aCPuDyVK7asaHhlSKLKr3RjEtmq8U1owW7lBHbZt3apNk
I5RQItFZbn6XoQmY7J7FdrwIxPSXg4Qo5QDpz2tx/A1I8+IpYUmHcCbZEcYFVnZX
6qwH/FtxR/hT3jb3H2a+2ZRIZVP3/3L1Aft+mOZNXv6SAA3puWwAojk6ptAWjakL
M+IbUfiW2ByHhU1PrO4uUmTOLNNCXJ8CdNfDMT+L2QVYLf6TiyCNnKhqhtRrUW9Y
DIYPEMXwpiwhK/6nFvfkiLYcHjJxL8Jwa2MU7YlpLde8AewccQj9sjKqZ1wnDzTf
C4YAjIvIsEyTLqaNHARM9oa0bzU1ArCO7C2dPm7wNiSBmP+M9xH2k0ju4foaWBHr
3nYNl2aXSNgZ6QVcLup2ikK6GwIBccl2UpN0DRE7CnMUMvo8i2Cq/zhYSjCvWZUJ
f11MWgvjl3A+myhcxDNSJ08s3r435+0MR/YcAnwjjisz+iaqHX5KMrlUqwUCcDXk
lwgWyjBiFrxmF+Ztvj0qXBoklTd5j8VtNdaHTfhXRfDJeYRS8KXQ/Q7AivfYRyD8
2MNkoSrICle/H8/t5IZiL/pTFPX7l+VxbmkZXrZ7ZzUGvr88qit0oIJeCXLbHQFs
D6wCVQfwsHBAC0iAzaozxhsmEZwhGE49Bm8BSBO5Vr5NDvvN8RIPx2yYA0MxIrku
qXsLTDjYejv2gNbek2qRaOAdoOln+zuRxWxEnaUgSQeI0owjxG3L1er3L/ck8Axu
l2gWvPdWAt3OtqxuYi3LP3QSeKLfZAxoA2WXmDVWEDOoKYofskMHgy+8gQ8bZTBC
tLxw24R33QbHzDk1WRPCAkQT+Y9WGMe9AWDbC8Dkx3GDYG9eQxn18DGTaKjBFebs
WuB5OCejXTAbNB+7/DmS+XKTQLsUuQoG9idSXjuCXFkhT13WzsmY0Y16FOSgJxTi
wxpkiPvjo8POo2QeQle67FeV5eKQIy7EkdGNTo7RJY378sky/m60cfpTE27+ab4R
OQtftTpZ6cw3pmy94Q4wdizwBHz2/iTTfU350fDVfUH4/thLzTQFGCT/7VSLbqTB
HSLRIodGbuFf/9bGUKtzEYMUGuLJMXGHT3qHuiYlL3xxBF4I4x3HS9Nfd8oJqCvM
7Ixk8mdGEMnrB4D+wjv/OcRlCddu4yvGxFn6oHX/X2xJ6w3QQf42Cf4KfKH01yzF
S3mJLQE/Ngd1UMw8H5/ck5PNwh7Q/9qXlJJzBW7jQXGOurla48rLM3Vcj8or2rft
r6xvf3IN0SeMHm9u54aCnfR2/ZWkMmQdIC2ohEyg2ufiiMi+EAbgk2+vCwmF7nGW
mO2Zh44rQ0H4g5MHgYdvDUFRBg2N9tdL+RHUkhV33JJPrblywQwm8F3ddtsHFFH6
gld6fpGSQ9ntiO7jX2iQXWzOEIq14tt96TofwHZfN112BDACLNN5dlwL1t3asiiA
Pdm1Kx9HbOytjoEuBrCb2J2Fu6w/pWJbeFVGVXjU5ApA3ozI4orL4P0u3HdepG0z
W+uRBzS+zhZFTsz235/u2ldx92LHfeUGlBiJzq9fOE5nrjA2c8ulYT1cOekPCztQ
KBCKAzq3SgpEiIa3ikawL33D8IlBcHpAeeHUYqoYawJ1Kj6EfBLibYUOSwahiKsd
EfE2VFWAjKsbdj8JN64fVFFukCkOUAgx6BMO8jOoxk56DV7DH0yEhjKa6Crc/lRf
uU/ThQNX5FYSNIq1oy6WguAR9IY1VYuKh3Q4REazdixO8Pk/hr81SMMAjkTayA+J
1V4Y0VJ5Kt91TwEj8GVLQuPaTyHm3Lwq1je/A1bQ0cuQhTf0tsCw6f7H1kUPLbL9
R6IEOwbejyB/RnSmUr5A5E5tRVIox4+NC6fQNqzKNIKdnCPbYZylJXTMrWoS0Nti
74a0LzDRHfkxYmdc3kChUZbqr4S46lb/i1VPFLeT1l2JC4YhoYsnmAO5hx3c7XsI
WT6dJyzF6+X5Mmr3+t4KMi17h83U+I3zAJ+aO6PYtiqWRTCYerDFA7hIedmuRPAp
FvLuyq49pMg+9ku+ZEURD6Wdf/V6+owrbK82qNHuFtqfpPHXByDorBmEK57apIuO
E8cWEAaS3SVOnFAMd4qWD51/M4daCA6XAK/JhK8oWBVKaQc1FwmYGvBEBwF/Xlwx
30S9J295Y4DggXcJ9pgGm+Oza1jqGoKGKh+vSn2ez9rrSfzt6RiB4zPtkbpqPBZE
vu+kAFxK+qrrBlB71p85Uj542n0JyYcQKUQtaWgvyBHrNA+xi6fVpZTZQBglF6wj
qguEgtNcgG8n7aC2Vgp1pMvIbNrreq9iDSqEEvqxDFwhvwaGZtG8SREYUF6+1y6E
p8ITJXK+JSZVGgSfdFem35ekn63cpckz24s4L9brmrkFXHgxkcBqMkgBMtO4sbIe
SnyqffIzBFx8dHnaNKTAa9IDDqeLMHgmHR96crajbgGwvlaQxVqUFY3wqw1Uh7Fl
hjtLNRLeYVb61U47Tv77p7NMoaK3B8U2riur5HGJsLJ/AcGoNzQAwHSMD8ETdUmK
Lkc1bxaUASGKAVf6Pr2KlAW3NJB97DonfIDT7/IMubU3MiGmu3wqqi54VSeOHTJ2
krq5QjzVHO6eh+btlDL547UyfqQQrzQRaQRaD0vMbdT1wLi1kgcbIdIEddqFFRmo
SLQbhMAhLIVtGmsBpbH8/cG8PcOZjfgAzhPgABLqid6BUSpGVjMBY2I67ElBU3jv
F6fN1Og3BhlHlVAjUphJ6czVLU6B/1IdoxX9nT34W8dIQz3PT6JMJRdXowNRiDEG
v3NrYnozIYpV36T700xzhLFJzdhYsKKHMZiP6hSpcCl5k58ONjH5ykLXFtASQg37
sqm6Lys8OIfxL6p2ya7m3h9ga2SyS0FvVseBllUDP3/xN7eZnyeYh6Nu2ruIqSHN
OMwgRqpCABuJQ9qkTeVQN0mupIZud9RvyOponNP5NNjo/W9gOZ+Vo+cMDdt1yUyX
qVvJcRMxQPzpNROFXiu1siDBVDlaugX5SWBzEjUEWmYttQQT7XJ2dy6HOZzvn2hN
1ZmnFe41i2XdSCBpthZ8+S6tckkr/sT2/YBHm67FNcIsyX89QjsHtOiQmMXLnU5E
tHpUuxRPpifFzkd6oNAnHO+DCHVVq19DZFyuh38eWRy2so8gild3Gu3F+5jO5cCY
WgtJTSvaTkuU45vs50Kap5ISWsLot60gNLrXl5fTeBxtjUubcS4cwmA4nJBT8wgW
P0lU5FplIeTh5GfmsFlc23D8U7W6D2ccWLDO69Ypm9SmyhDmLnsnPq58CIQV86Hd
Lukus9efZmucKxCOw7ItWiGltmPnLOTwmkP8tVn7jz53GP/YG9Ez97FDDBSpAtob
voz7Y2tW0l+dSLUkupjcj/CL4FES907Vl9s+osMuBQRWlgkO1Z8L3Q7jGcHFPKm8
Zbut/pOX54uZKMXOn84cDdhhwZP7ns+wvU4BtqQY5OT7zRbeh9mZywBrL4xLTTVk
9c+nydYRxtT09k0Trc+rfsxmEbehtTWBCz3vKRExoMKnXgQn9O/EHriLeh25qZEl
fj6cYdYHx6JI2BaX+rYE1jPGa0koV4GuwtRqkC5q2xzI8Ia9nI7UhGLZ3Q5v9VKD
m5wu9X8Thx8D6TkrfrZ2Xg/K/U5/wlquWpGWkUgxBSErUqfxoTw0wc1gNJoVodsL
48i8jtpFjSwBxy6Y3HYC31kYGR/v1b/4egj1og2MG7ZEMIlJ0D9Pi+dEVnzwRcLB
lTvIBQOcxavPGVfFzYlfv+PKmiLP7mLC2xpTF7KtMjJB7csQRGgtaAK4M2jYqewg
X5WTpPNlImS2k6/OVgxUUHjxjHxMYaJtZLuxnAnEoLDIVHVyiHi4Gcjh8FvOjtIb
3UlNNmcdtnyOfHLF9krp5Aqf5jzQZBAvh4QzBnoZx5Fax5mLOVtj81o0CFSDz3Hm
XidWKdxBPZrqSHCjofUlGldw/oKoY7zOZ25rhVhOUfAs8MvTJ8AneVtaibf5kcPH
lquQT6qSKgugMjISAeQkp0qp7dqPe/11/6uWp4Ex7j8ZSLWNYeedJYByssFpZvuj
vUgZBfCLe72pYTxM8SzKul5yefHiNRSr4cT9ZKYSyMropDXMsuJcMW5N57AQmM3f
gUtjxhNc0BUbAax7VLcMe/7liUxFlEColMbOiyCyL4WyfMVmyDGn/03kTdsx5SVs
Qe2AQkiE6Mriv0hSoRZ8znX0Z1p0UV0xg/wv/ClNsFNl269EGop0VmNINMxXHezq
KEtRnPPUoiJja5UDn5I6Ocj9MRvdmnrSLi2m04GrPSiYdzNyKBeqpTFa27Mf51W1
j1ThqMwupRAl0iLOu2Kof0Lh2nWIB4LNkAd8BoGzfaKw/Voj8FaELsB0vKKINokF
UUCa2KpW/i4rxa6E5xCbBo/gL1pj+vrce6AXWL/mvbbXybvwRt0aehWNACiP9v6G
OpR+YDOnF0iDSYTG2BDOysWMrPcuN2s0Wi4XkMpc1No+HAnrHR16QA9/pzXoMlaq
5/1CX4ffxoD5XG+KVQj1cbSa27bh4j2HjkzpwCcsXpG4TCKNsMTnnv12fjfAd8PM
OoHOR2aeMxxlpCMesfnKA+Kt7rSMrKbcX8bKZlgjfYr1bYUNwrNWR23mPc5G3Ol3
+g/7J/T3i7Mll09syHb1t4+a26FF7tzP41MOmgvXVR8dea5217ICktwDhtW+nmKK
1r28kW71eFSZGmjhyC4FhbUrDbEsQyLbEWrF04ecI9sb6eJsSzEpxKIzbPFGxgt2
8qqxZJ5PrmQHjHDcx3PLAnijK/7UNTDeLcGmGS12z+u6RokkuNkMB+uVRxgjBzdY
+CEldIj1k2a+13e1exNrdonsJDM6Yrg23OoAXRSBVG+epQKNp4dEMTe9w7z6Zv9m
Uur0kGSH9rXygWoOF8e5/c5iCpBXq/fsyLAkudBPvaRN9JtbhyC+3DflxYRKbuax
igMHXwh9CbZS5XyIgZ0GvnHLUJD4xXCOaViHRiMVPg/ExmBQmmmgG3W8AgZ3aovL
YJoPNgSi7F53f+HmJ3TAAtClbLC4wgUWg5DtReWLIacdCIBgsn2Zq8E6d4HJSYGN
p9fuonZgFWTWjKQ5iRSRcP2VtL4LYhHqqVTNWEQj4FiIEalDrkukestk5UGOKJV6
3Nq+u+nzidL786BwviNnfEpfSypr9hgRio6ty1BCjd6BAI77c2Ma/dNbMTmitgGR
DzTPEpZTp3obmtPVyNVb8sXDu+/fEd2lPWfE7MDCx7oi+jteQKjOME3GwY98wpnD
2rz4jKUX3dT3gV94p+IbiH6cGLSWerQewQD+CtsdjxDqsZPjrzrDlGSzMefqNr0G
18Y52b2ldMDbytGVy1TXNjvRUssLCy3ho1nc7OxdM3/7BHICWupBeS6JfZ2mOBe7
GWN3YHRTFWC5QYJz5a7yM200cNhU0bfy9Z0wn+1K8ePP/G6ir/3/AG4GVXdFsHGh
Qh76MxtNtmT1tx1+LVb1aYdBtQv96T0g8t9LCn0/yJC+bvnAE+zdPCRd75udWgtM
Ajxs5GMaWs4uUYxY5+k+1KNkhdry9fLGvdnAc8BKvzRHV6/rwcVom23qoGvMRwYI
h3Gx7TUs8Fhjy9BZbiCVKY0aVtn4wNDomaQ2Jxbc9aAeu6pAL3APiKx4o5es4M8i
O2ydCOmtGq8UCk+O2cRhl2NcC1e8pxiqq9R7feYhN83o9TJfo6CZiLiUqo/eyHeH
ng3LeIFpybr4AHc+qcae6TxxSHrWA/H9FzIHBKE9YYFoulmYFH5SYRFc2nqu1vid
dKeVoLRMUp6RBDG2qcII9AUKjyQwisyQOozzgXhBqb26Rpk2cfJhXs6721jQxI0r
HvQwFVQEmU+xEZY+EBbdakqSfj37SYYAhG6SCeOSS9vwttjvnX/1KqL66xfrsKd3
YR923zCLESmOpNr04XL1qnxLB2P5HFABZCO34WcZdwEgfBFSv/gbYEnBHnpoZOta
EUQ592OmWQXJESt3bkv4WeAAiMtG4xRaW1PuxJhILnadWVOWxTAosWzwDmF6W6sO
HO4jE/v48BjHVBdyPnSN/+yh4GNETFnfg58wPWPp29HjxpiOG0uFYN/k7gRYUS+6
5AITOBY/iH63CpfIixHT4urVjDFF0YSGcuEcICx2pc9KVqLDbdoFdONsCSUXvqIW
obwnV/yRKch7cmb56U1ClmDWBayd6QPaNjpnsfrQ7r//TCsyxr845OjJ900BY3/3
3ZZH4gWcSH/G9ZN7SvPDM7AEeiONIIf0tJDgxIbiCnj596PCqAP+0aQae6vkbmvo
ZSTDWDz+kVrS5cKLapRst1ow+Cs+OjKlDwV23cp9tUn2Lg+1P+/j9BiI+leZxVkT
OjTpaKQmOccrDHlHSQ9EjRWtugEKcC++PPF6/LSC2rmqFA1wenHNpCCYADeHCIRx
ueUC2+tmVbQmUuqdX1Zaw10rRmODEISr4UCLgPuwR5iiAD1mkqO3S+yg7LIlFJY5
p2szdbBUPTeik/BH0mwGvNvd4VrGXRMmtc1Uw9fuucI=
`pragma protect end_protected

`endif // `ifndef _VSLIB_SV_


