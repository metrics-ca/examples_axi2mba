//----------------------------------------------------------------------
/**
 * @file vsl_reg.sv
 * @brief Defines VSL register class.
 *
 * This file contains the following VSL register related classes.
 * - VSL register class
 */
/*
 * Copyright (C) 2007-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_REG_SV_
`define _VSL_REG_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
CQVKEuFVJ5/zELlfgw38hcToYaEwAyhpiK7gwk7z6Ap2EhsHXwEdfb4xXIWqs+wx
tIQKhbg8qo/UREgUWivWjf3fiSbQ9GZw843Pte8TxmrdT5UPQxHu8+5e/kG7OGku
guL1a5LO2x9REdvlGA0NAk/H5M/bG9haqk6aSqYxgIt+BYFAamgPFdpn/yN+vZVb
TwlyaRD7zesOvGXOIhPYW8tDikf/6ZUX6XOR1FpGWIpHhlb5GdbUb7h6NB+lENsr
4GMEUHf/xgKa7p3zErl4JPsluZ7Sj29Cdnw3VV2+fQ1uMevzctorsPmwn5eR6H/6
EHIHMhquiT4VApVEk2eQAA==
`pragma protect data_block
1W63LBKehqsA97mazU8ifTGkDpRX5mWQYoROBnbBnuD47B1chQNRgLBq9J7j6SXM
TFzg93p9cHEsLmgrMq0X3zp9z1r77hkFlYc/fYVfQ2jP6XYbdvBIsoF24Mm/0s1u
3bxj5W3kaEs2V5IyOtV+zHnsVCcOg3LvKEZemZX7AMXfhgB5sg9eDnFRnvzL16dF
jMlvLJb1fhDgksZb2UzA4wxonBcgVD7NnSpauEcSSZE/qTsLdWi/5/ypWPxQkPcA
K48o1ifxnn/qTWClTDwdNHNMFUX8w237IXfaHyaEWV7rPuPjtQ9sVLsLy3INc9Je
s7P+9mwmVSWqgLICLLiGhLrW7PBwpikcIG3Jty6kNqnCXc+HmEssj80XdWbCWKGT
0ORmlZiDrRkYMNcgt5qhmGkxpnhjzef7swTdO4aXBoQW0jG3szEETQYAVgRVgjB1
r+PK9sebMN0DA6fNOynqJk+6XcyoxHEt6OMOHsXkZ+QVvezHUueMtSGOW6Hm7jM0
NQ3VAkOUKU8GK+kjQ1f0y6LuBEL79ADG1nBvUb/hztUI7g2uxM6pnzH4C4ZbG1fo
nDti1XsY5gMZO+3GMiztzcl1iqOwcG3PlW7UYJKYvAFk9TmF05NyvZ38/W5j3M+Q
2lVVm7CNij23Gi4sk1Do2rowJijkJrVjIudYn0XbZzF1HoFU66Evvs3RusCHSoBQ
z2+Ol5l+VEoRs0MovW7RqTLufMdsAlb46M9GGVYJWKxMWaQW5hJuBYMjOqf0JEwY
3jTFDAQEHA6Tldo9P3YjKgOLTCPxYnjODxjSUVbEBTH2NS/9ZKCvgh3FvQfyx9dI
dyu0Jg5BRp7Yd8xuxtAbcEV1Kidq6v8DQFSG53fFAdlwUeXy7r7Zl9JQqAwf5lxM
pwnb9IlPuWLyC+FwtsnPi14/uTyUZSe/Uy/LAScQ4gNmvFh3/oCNaBOCKsZP7763
8SsWxhyQ779+TxINx1ayXNGBPmNlr6SzxExz80Av4L0IcUp0tzV9HB6RHSDUkdnX
nlOiz/5U/BEc/smEipolbOLDElE2xqRp9ws9bR56xxAjLnmgcdf0kO0LC7pvDjP6
7sOeMSZcvbKx35IF8VfXO+YvAz6steFDwbNpjO3HMGVX9oKC08F/rmaolY2HDoWe
KgcLEAqm6SxhqB+nJ5q6XItQwq7x8o3XH49XB7cCAIPJgWGxbAhYw+CS63cPx6ta
gEtpiLP+Ky24NMNMG8Xt5LVMv8cc2Oh4ontwVnEHhfCM+zJBV10Cj+0x3iK4PVaD
E/baKi4XhWsTE1+OXEIF3iwpuq4rHAergDHouFIIO+ZoboNj3pNkulTIzcGkX/GB
Shlwozj4ISN42vv6WzhVte5FuKF6tpwliZHBRkCkwknel7gZdqXfSR3t5emqou8c
CN1PpOf5nkyZu9PChi/Uik0ScnGFwMIssdGGdiYwVcJMBrMyNyNK5fS+uP4rgBq+
jrxIhjKz1iP7ywCm5vNGVBMkMwRejDpVYdKms0g6cdLrPsBvWP5kNFxIscEljxeg
riMaMMfwpwiU67k3hm87WL9hMe+6CDKVBirKZlrzbI11ixJTDe0fcjo+2KshpCnp
/YStP4/afn0vLXYPpofes6ePTMm/AVfHkj4HVF2kEuA/XGgjwBLR6V6ypzjkM8KQ
lYgljbI1IwYM60PnX8Ds9HgpyWkKkWjMkUaFrJtue5Liirp40jr2yVDpea0rF4DF
hGoa/ryAdQxK9JVBeJUyC5T8jD+BUnNW083pY908U7GNb2q/Sc8pWcM/i0fObgyR
G/QtYtTs7ZMuHYc6TiBz+8Zt2TjiziWuL3UAIGOXl7Ez9u2lBRkGd1Y+lW9LgpAY
ZR/N5dSguPPXD8Is7ktjdP9cP2eHrWwvjWQiMl0EthXiLq2EH70FHwlTbTRtcWNm
xRxh6BN8gk6YKpfGffD+/qLknLg4vcqdF7Y5sth91PlUD6hF3S6FL38ZVMo5w1eP
SdjQirCVJ5G60ik8kPpcQV2l7Wz0+xFiM97qEvDD6ZyEgFEH1Rlh8U9TohudzOlL
a59KwGLSvSpQrhOfu3bqhlZ10Kf26krIjpB6R9EdSUubrfzA09q7R7w+VHwHdann
QWNcg/BgyqrBRvc1YbwrltwVckVsd7fsmGN/iiCXIfYXMretoOV3tTJI2V1knhsR
kpCj2ohez6PVyAQ5o23723Ejb2sYonBxbIIJuRL4Ha5Is+NY0LF3B1d+Bwi0a7r0
K4MebcjQ+Vic5OSx24ZH4OIbZQX1kFeMTHf4MeZEJS8ZP+JytD9XjpJaApOGvD6S
pLHIIJHXJPURWHuvOQv0BY9+8wb9p9h0nbNydhCgnr3NweGx/2TZRL3QchPGAKVh
hbUjNmPIzL001Z8ZGmgWh3126O+v5HcyuJEoaWk5iXkk2jTNJPjj56x3J1JNBBe7
obb175XUCUdl+zqMNewelvK3cdf+d+flhH5numyrv+CUYiY8h/6yH9BrSpv9SdgG
0CLTs8l24wJqzXutLrmSaPPd4WwmmFPRr/u62X3WceyFiT74g9w7tffxCC3DY0pR
fKG8BPivh+aOUjVexfZAPCHrRlwAVNgSBFrukO1wMmwj8iU9m+8SIWbF5SlxQskJ
ajGkCc9Tx2tCVsSp9Q2knIwJHHEeLWwJcpwmq+liQZYJQPTJX6qn1CYTzCScXpJk
vJsPnJYdAM/dCO1LA8sLy0TjNFtSRh/8gtr5RWWBeSdq6ZJMqtjiCPcHEV92IqYt
sBXFUOP8W+EXe6hCXeepgG2endFZTRomdn33odTDrXSDiC/Hr1Oa5pgEcctVk6xn
XLTo5HHAUnkttqDL4WqCZpsFFpJndOFo4AbnYnTvPNtZXSqBGSY6rtOyJ86tHKTU
v6D2TPSigy2UqI9nMAxCZW0VB573leW8MCMUlyvw9PyUL5Hv/wOwTkzDjx/Rj+zm
U/OuuzoRiAP5gKLviibj2vjQEbHqcIhYkbNHwe6xAbO6rur9hB81/NEW793+pelV
2kX9b7PAnNnUCEs2Qnmt1LhBNTlTVVZ1b9LAzKnpcqq2ENBtUcNU8DiHYFvZlMA2
79iOIH300bS1t/YTg02wapZrqSIQBMxW+4RwjzFPQoCTSSS+imnxeFjOU40Isz6O
c2KTb13bShl5viv5xJn/TSy22ad1jM8OBKXnq197Q1yIV39YcrUcIhs+og/hqvcU
nA++3UNxYmzxnaAUCtGTgtATwwpez+JJuEy1DlEAN1jDxDXWVZw19D5afZgQBCCS
e7BatNFegtOmpMa8uqSfoXKGCUjBsovyLggG8I7TruZehHKa55SM0wsUWhZyk2+z
87LwyX46J55VPvK+5Z2gN5pV0zANWP4mBNY07TuFharIXarFKl4ML4L/S8FzhbFz
W5lszqbImninWwcFbgmDn4C1HW/DAK4FzyMS8Oll5ztkz7J3NjrUis2l3jjd/q3S
6Qv5TxRQiRWtoz1PsU7V5CWVd+IzxuYX8oHVA+4ldu5S4r0rhQlxXhVOttJOGmc3
n8tUV/YikcW6lbUaPgBo1qzXBpPBGs3nh2FDj+KBDBLROxChQ2NmwflILnlTJlbV
4qrEU7lxqpvhdWzdYosdGOpsTHF/4NbR1NrVwsoy/g33lhOYRFkk8ANSEb28j9bK
SnHJFa8fSxlMlxZyNCueOs0+IKmdzlAx5V0sdHIN+fMeFNQGXDZSRMg3APxhYhuk
GUH3K4p42pR5Y5Fdrj3SH1AjkCTeMgoSri07byCfPVX4IqIq9UbD+JzJbg0oZ5HP
yffIk2VpGydtIPJoBoU4SA+EfO/w58loW1zqFc0HqA0SIJIu05rF6HZ+nBmU173R
W95WyvS70KPFdUH0kzk3hgd0JZIAdAesILSyHr/SmwfekzfLhup3ZIsGqBO6IZkg
7orLFPIQfIME3DQTaXcyc3u/k6To7Vx9GzeFYb8BDy2vGVIhYKvu98QCoNTf0gMU
TXH5bs/VQ0erTiLk7EucINDzwtcdM1HEXRtikPQTHGol1tQnEy1+e89X5qRFjRDr
kcI7ci9BXbOz/9h3uEXPoGNS8T/gMTpYjNGYPJL3tUhMxoqI/dL5ZAHEf1Qfw5yj
s5Wjh9atcSm2UT38JXkIKCcRrSG0CBpYCp4mTHQscoDNJOnkeptGqxmuatJ1Sl3e
2aE6bwYxQW6tIWp7xsefbHxKTTrjjIJB9YlN4bJ6w6a/jKiLgJ+fOqvIKa6dH1gl
/dyF/FTpVjZzftRU6NWQT7xPmMu6spZYRbyF9gZnf4g9LYHkSMuhkEBU3pMC3GP9
zrPgL3Q5AH2i8ld87RGjafU6KrPaiMQKFkJwGQNpaDKxllrwA0UQLz1QyEL/3hVB
vFdOppyTc73w4jCU0IWkwilwT8CUVePgw6ubLWnptkbV/4VBeQqqnTvJ1hkWG36Y
rNwdob96hmVSsPd+z6N/l9LQSKvWyGrFvKAEqsPu8Lg6mQAvOoCNBnye2wHCSkEX
7XGQGKsm+egYNup5EnO/CNyDJ7fQOYOAhS9b9aRY63FP/7TsYHxIJgOPml9+JHry
iZK5i3rOy1vsMshitI8Z/gapZx5pfsnaiYxC8IZI7oQV4mcEyyyPm/Lt7pRGkvus
ajP/6YVGSkpwOvG7boZUxibKRN+GbWIluvULedSvErB8si8cnhgASH63mW6jwrvJ
5DQrlNglXVTo3z/WMD5h5On2q3A1lfsCufX0GOrvQPAmlHd0GPGXzcBJasunBe7r
wRtoQ5gUJlPmGgliUqvRb/2a7Qo18/vkX2dweyf6PMhG/WvsA3f3ctjD052TDObW
M92RKAB0OcwbgBkyWPq/4GX6X2VLw4St1z38OtaoX3N0jj2+6txZ2bVNM3gUVftj
UL8GNfA3UB5Usv40cGC1RqAZzdw3nQrkeCAbhSse1xxu+3Dli98KjGm/BvaDupda
W95+2qO2vDPf28dvsP/2CYFUlutgnXAoAu6fIHx+/mLjRgLcgQjNYn0OvGJI4Gmc
7/zx3hhN/PRWH+FhleQVozX4KKKwIe11Bnvcf5uDYF1y/PLck32OhbT6bMyj4Qvi
IZvYtlexn7+RFS7oeQsR/PfEK73W8PJCBA7l2ysNtRr/yLT/nYRWhubcTErBZO0c
+r2hhw3TDCu9/P3VAk8ZOtCBVrqxbe36lvRbqplnD09SizUh7Fp8MN5LzuExj27F
X99vsOvUYwux8Z9NdeOLTYqy1PdzpbVyS7YA2PDy/BGko6JdOlofemreIHUAQPnT
oDBfF63/KDaG2BqmPaaKPTQl2+Fot8qg7INsNePpMFsMPIikJH1EKCETxr8+xAqq
4+ikfrAV1ml3fC1dGihnchj7J+zd22/HOO4PHGvnZPGRKsCnR7BUMckZ1ONE6gqk
yjX9vn+2OczvQ3Rf7g34lGL2E3AS8E4XbGM605NyA6BUxn7P3ezHwyJR5XLDVec4
63Wm+CNFJkvfssdcshbpXHszAKOl8DKJHuABZVnn4cQ9NtKtRz4CgidQ1DJ2r5Ar
vRaoe6ZuN2PlWaEchmjeDGevzh56losqajsE8WSUfrqUrLXeOdaZrWtznLZM29fZ
Jw13HzETyDGYg2ggJPXU0f9Y/TeIbSAMAEYrt4y8o0EpAwVyIO5BD0TDkWFDUJiH
4ht3sr3PjKyFacEyKAIyRFSJ9k5yhsQvx6hfOCjx6DMjBfPbf0T5BjfvJWgG+KVf
xwTVVSoqEKzTijiOuU3DEUM6+epeLMhyWed6+bnTImp4K2qaDhTWayihktuBmQYr
YPXPWHg43cv3+m5VLt/kzPN3Qhh4a1p2OaHjIyyiUWIbbCUQTkpYcOzTuyOWaNNE
/PIeOE4RWBhgUYtypji28CoMT6JA1jv3e5WSBORc30ox2gXms3zLrIC3CTKFDnMo
TQWVJBkaMXbQgmLq1NcI/G88vl0PhB4jBbyoEQSVopyxJKxpKvC1WrnLv4SHL3dn
0nQmdCkMc9f6EKuB+o5wL27BucHUKkN0NsfxYxPpFtXfMnMgLR/Z7SUY0nzZD2zn
MxHubElEU8yFQSZcXLxoHnI/96TDuaUuHHeeEdwOZYu5NMc3cA/zlAUKsRMAil2O
t52GtqBpHP9DGM0fmtq0fFbg/NSNUWjWrINtmgEcrMAqTCTbdNmWFGLrYaxjxdVM
hkbe0FZnRw5G/FKvvFK9DFGrKzWnTXHeBCqxjs92wkxZtMlkFQ2jhkQNvN8j3ILl
mgAfDQVZenpPK4Dxe9V6XsIq+4V1TkwrmNlE06sj9OTEX7mkcZTApag1wstOkIVJ
tzgq3iepIfZb+Zr5tpbUkAWPevzMIJ4BMcnXjK46I5FTyEsZOgTQlG/V8cQmJCEd
QP1xsqrbMPKpiDg3ohsaxeEfaZZpwl8lpEkRC2N2AAHsdAocPLb1/NGqpeGIkeKx
oHIEz70ab5j8y2OlNvvHsOkOzQCBo530nswDcQ6lZCARLGGh8MgY16FhI3wVah2r
OsQl1yROSNokGgx6svtr8yrH0kMC8oFzA2f4UgD3/3f/fGGIaJ5Nk0HZHHJoNV+3
BQuAk9Ew9Pebnb/oRBFbaYOvlVUe6Rc3v1jFUHpG65zaqq8LkGJGefCi8YdN7lW5
X1NC3kJ/X57V9lk4wxtDVKm4mWCsCPStjUqN+vDkNJquikh9Wj6KwF+FMReW05GV
rIyTbM58bpcFUra4CcGnorFwPfeh+QpnuH38lUG5jWKJ4j75WAztqdohTihcskcv
oX8xw2nEm8dTVkVr9S9/oP6N9fgsWJ9Dh6MZx0WgvC7oXWlU1qMC0QXQTP/F5YMB
etfnUxLFMHbHYOVxpNt9HpVsSOSAnvBdeinKrbJ5r8HnElLlWcJNLJzpqO+xyyRU
uj3SmKP6b5/YTSSwESiCAyjVeO2dPsKjQsLenro1oiu873l+HVplNBMQPQhHi6QY
umIYlVG1j0xYA1IizuwgF4FE41tv4VAVLLE3ozHcMO7QS2HkyvyWsVYzQPZph4A4
jmUoZiVGEoo6IlY16A2ta0BKa8giiCyrcCoU4qZd/qVTeWcpIGbQxJgdZ1fI6DUD
4IkE2X3/MNj77REZxB9IX+52LsS/nA0VBmGUsGJfsYyBIkc21pbdiiUp8aUlqDDp
Wj9bE7m5yNRg95mld3WqXH8oCkPluW8vnR35k+Jl9RAl34evXhBTt0xfwumJ1CQ1
dJdcO26pC86RLeZhjVls1+jg3GNYQHwJsi1F2k+q9kK+KB9vTRY0QRqV1AJ0etb0
rKb2EVUOslVULNaGjfi/INsBU3z8wEd5kM6i40XRtuQFOTocgclilGgs5uX7kJlh
cI9nCdSqIfIHnJi7tNp6GWxa8tv2B1Tf68YdYHvQbbiMbyc2cFOBRTT8WuVzvbBb
PLK/RVF15eEoKWsdma/Aa8p2wjHk+K+Xw/GReugRAQgzkoASqupm3EXrt7BB7owk
THke1bt+X0ibcEF0oeGQ3TSp5+sWj4SYyUZ63fTH+wcgT/fgrGX1YRaRjWRUaxur
D9SkxbxY3FA3Db/sKAJdHiVwaMsR6CcKPo2GMQOFx3gwLvXEDQtUcsMH4Uyqg8bb
VKYUWoQVVF+9f1BS7IE6Twiax041eGH4XjlBH5y82Knjb/uhxwnC1296dNyjdJ++
oHdYXhl3/cQtztd/Sk8PHxMpJJh77sSwb6oSuGn1EPsL5sQTYxjrN8R7KFpHW/rC
TRkFhgRvyYQwm/879u4mjWemp1loDStY9anh+0yxfFZrohR1BUpLgBQ87nlPBKGU
+DjRkCcQuTZhiCpoYTet4Ddf3C59Vz/x1JS6qARrh2rnGBOriSS2XhoBTpvIrCnc
ya2B6hvOMRYgAv5AsPJiNcWqDLr9IIGhMdD0VAqknvM87KRrx2Lku6bgIfePWgd/
mVBPk6CsrPi62a/vH4zJFpbAiOf2F0SlT3/Yf0zj06ifWD5yDHdhb622BzpMPrvC
X5e4H+Z2jlRHeGBYYNc1Li3Ue9CAx4Ldu2i9fEayo4Lq4ZSGabxUKQBTkwxOX1OG
/574j0VNPbq2y4Nnqmvk2Tc9j4Bplabv/qHZnQlG7QtoIDDBZnQ3Lif6aPFpd/G+
4Oh8PRblwg/N/xou/PRJ2ijHmA5bLwSDUKfTYEIEl4+8j+YzCRImF4wUEvA9TdxL
JcYQmvRL+gtdQi4ZJiONBaHpaMqJNnWfnrr1XZFuzRlSwoEsofGkB8kPDypWTeFx
77KkFTYyJQomHBRl0SlVqIul6AdE815gI1lnspDs6RyhYdkoptlYphzwPHdrTczs
Hq1h6sdMv8fSYFygFDb//7AjAORC6jtNGTCtKNH9ljSaLZT/LLohxniOylGfYEtt
OWoA2Tm4q4RLgjnltFzRr0Q1uO3tNw7/rkrJ1xDxUfaNqbYBOo/hQQ5OoTMQps6n
hfIcpQuPQNFVN7F3wu5IM+Soj+/JRq/d+vMEpk+sOrSJLv4KfUtP8//RhtNNnFTb
3K0BvElcu+JfnXT7X1eBo0LniSxSitgWE3XxQzeL8cPZB5BFMTgLLq3UIh+XR9ok
rPss3eSea8Aqs0oo7gQOFHRoFZ1/YG88RVbdO8le/zF1GCQXAZ5SC+3oZz8zttHd
PWnucO2k2TMCF9JLRE8RHi40uxAnaMe9iP7fOJGOVHvFHzT9Ci3XHqZqPuxZXbBB
+jIgXYmzMYaMWvr+Uheowm9PEqVx8B3KyPltYyn6bWz8IhLlmmLsPmwY3Mg2Firw
M6nAObxVsdIiuI0i3zAsXQ4IiXljWiVaZqJ7diZSRbghJKYzQvplzWMH8CL1cayI
VpAHO3+ouJg+0l1HSec8ooJE7uwKCYNY/ndeK1d5w9X8b6XZA3DATt5ynL8U91wb
nk36it7Arkfd2kZrh0LCwPg2ng74ehyqi0nmY+HBEVhkhaBv//OoxfAPwse1GQHS
SfAARDo3j/lX/eVFNa8F/JEnflK4aqvfn5au10sg4WOTnlXfYkMzOKoQ8oI44Cmw
2Wo3aB+VkkOtD2/5rKJI51E6jSkY1ft0L9JibrBKbKl7RSeKkec3ynANDJUp3TFQ
iYRxNnA72O4dtGK5vi019bzslfWOvQQV2IdwemX05g4P/h0orbWwIEFBImA67Jdp
aDPFjZ0/+Q5/N4rI0+AvT+xiFfkrdX+C0UWQln52AgCmr8UDbSZJcRgRtwfAMf0g
Ssy8WnYUbglLUrQStFjZWvklzPMJvoKNReZMO0wOdCka+bCyBz/P+8kBhaqJcX5n
0Z9VSmVzpm7VcU76DyMDY+qH899NTbjJ9lAVWpK/mojZOGHcWAMUJO0k1W2n3QgH
wi1/6IwrCdv283TK5+hXYchjyEAOZH1muJV8Ts+VcXS+oIdjj/7S/Q/IyEql10Yq
JiaiwHJtXHVDY7FCTzQRaunixaDmocY0VMNthcE7PwkXVIVuTzGVI5eB641/y/se
ZFmZuHIBEi6KXVn8qstb5yrOtRgQV50TV1SV8jJ0AAVnrWYYT3//rig02gP9Ktpm
yuUC40c/glz8W4/fuzyXfgsn4iBSB/PUXhIBuxdKF4KG91B1DAVWTZvnjUBfBzKk
nSbjexgES3yEePk3LKEQyJGOuNCTlCk8U2ev9GIHP1OrjsuaKtcNfkvEISKgjNEl
ODOKCH+5b5qVfPZByy0yhqelS8iPbtvEcAqhnvPKiNhPDavX+oaf1v5YElq2obgl
EfRnamieE6sRFDDVA3UqUfIVvEjltIQ8/0k4SajjDJGqBmhoBVU0fga4EcpLBv9q
e/ZLQ96QgMyzSg3gLPrZirFvqoCgaxSom2wpj/lQKgI/h7vxmcVUkWGuO77tWYUe
zIGRn6QZxXxHq2OXszdrOB1EhTkj9iaCa3MxktoFGN66T7JGvFgQxhYgoGDouHQL
Tj0pgLjYpz4P+grA2KD/+GBYuJaIidwgfZx1EdHjXGvzj6d8N+BGRe4k+/GSiOdr
IM4pfuPeBSOLPLzu+hJ5uxdaK/koYOIvGmBDCdOADhPUA5SehgowIp51PnAFO2lR
0Cu/GDhryGHO8KLTd4XSvk8d8z0DGl5dBvK/cOslvIm+TTcA0jGI8RcfxlEtGzke
GOXy3F90VEr/25Cj1iSweax3wwfx1bNUyBcIrV8HsSpOfhJ8EAb895bRUfhmeom6
kmRfcfaufhZz+b/PQvNaZFSXCLQv5XMwkwDnPkvfo2rjvGbKK6oSs+SpJdONDTpD
udX1r5Wf3vkqZptDAAOn+cbIKsrLy0MD51KVuH9MtsrNXGADtSuy17kdLyr8NBaU
PjIh3ikJBbU5Sa00plaLypRlPn/hKeftK+oAsC9s2xTSg8BXB47WYHr61sD9hq6m
dbHJJcoczvSCCKeknQ064XIvhXRYrFfgLs7Mw/FUL36hGhqI0rPSYyJD/Q5cdK7z
d8qU8Un/EnM5U5WjS/Ci4RqYbyRZ7COUtqapRlZatn5A4U+pYM2CWBy0gN23Z100
qpPRLGnlTu0tvl8Iod+Mr3l7FByb5E96yiGb4ATaW93QOVCsb9ha3BkgSHk38N56
tN3mDNnj2QNOMoSmg40TOSaiJZx0Q0FvgPhaEcXtb868aP3dvEqJHFAERQVs5bqB
QUWYEKWNukWEk3skEXywpujfQS4QxZNMpLv8tlPq28ImiXIGwryzZYB+TZ+F0KQM
urI2smzf/qNfeLh3mGXEnoOOGiZGGfA5YpyLpMJduBVP0s+/yUyQqWLOf3TMz5yt
eHfrdbSvO8bHgfGX2ubzIuYmdwtKE/F8+/Gh814BPnkPN/pXhcdXe81Gqwt9w5Oj
nbXGqBLiKnF6x8Jw7muhyaCQElZ6SSp5Fv7+nVdlavhVDBmXUYztimYoMixxBSNy
1fHeI3Zjk9HpV6oGfDK3xhf/dlbbeXgtr8KkRwrF5ux2HNa8iZITE7uX2k0OAcB/
laaBpzD4j/BjnoE1avx1PjuNF498btyZ3jIGT57sBs7oaZlvtV2pxqw/Qb1+f6wg
AWnJMYX3O0T9IbKIx2005md+MnDIX7h7xDiogI6a9dhhX1D22aOMmGkt/aYKhyte
5+RHhG0zM+OEe9tfpTZuxyqD+r5/qpDTbJlXU+RbGcYqrZZKHgq/hLenCYGOh/2Q
lJxnDUngz4EwykGVS3qh10boks6EBx0jQCe7mIStuP1eGdL592B/n9NrTLVeQ9tY
Kq3Bp4rA+dhGkifnTFp7OoWhdEXiF3S6NC0KbK1ye/CR5Wm+iSxQGbdtI7ZvkOB4
iEek6lpX+WdCgI6y/kNy+iyKAcB20bGHMatt3pgqcZmRubVfPnJp+OV10kpVtVHp
yevtFby92seM7pdNS1b0osDDzNDmJlvgiJOZpMT+qHQCzgnY/YOMizf1kbIvkAGG
nzfevOL3AvvQzSyhKSTlAkNtjs1YJK0JfoSXuTa7e+7NOr6mESz25MLCK7BTD4C+
Ba4vn+90N93/t/bQjqp7O/6a47OeeLz0mlvQ+Wx1Bb6Dy9FEfGgDxtZt3/7/c/d3
biav5YBeXd43UgpTbutjBkPrXeqJpUSDvObas2X28/h0qKWl0bHCHl29tXDdKjUd
qcTSsyGnU4TCCGHCmWQiUpOyvKvoxMQboveH+a+43Ff2rZfXwiFDRODnLupIK5oy
3wuOHX+vfcq0XRYYMy8PN1DcG4IlHQuawJpt3+fjFKIUidGzq1ZcdLOQcQhL9S7T
PiGspFDI537pHTsouPU68XVKWdLmGLzrWB2A8imAPA641ojp6fH/YDNTXsbED75f
ceUZm6fBFi/1J9eyBUk/zI4xelU6Mi+oY6tEoqr5spPWg7LHhGKNeIt+wRjGNrtR
2yQEk2yYMhAmVC1GaB/xGYQpJs1HGwQ94hCGUUVrS8g546Op4vjkE2hv+2tk3gZE
9O2OOJ8e2/Cf1ndfXZtTO6w34IsB5xzq7b6QmcTr1rRBj/TwQy0oRd9m/+rsWQFK
gUUvdPSwoOPtt8lHsjiZN0T1rEpMNnmKJvGem/ItOKKT76mbUywJJ2VwY8Q7Opj9
Ttdk50bSgKac0OUmdkN9AVWmxTr2RrM9w5E9Hz0LzPG/KZVgvpFSNSjx+v3VLJwO
tryXWGV8lnF/tweZIvX6i107MWr785SSGcW1EhMWdeVsu+oqTyJlzhxDJ9vVc1bR
NZrS01WvtA24k7Lr77X4o1noFnjWw8UFiZV9jsP/gRFxv3UHqL1h/Vzog6kD3wFw
mYIWVcOgyJczpwzlHll9/xVZ2khyMBRm+TLJVt7fTNC+7qG86Bvv5V/GcXUtuWIH
SHVMtiGFbQgszvGRvON0aUQPOqOi6M5epzjLkI2uI6alji3QDIwGeg3WKyvLjQ1C
ogJPmt5/Gx/rk/ztXJNz1sm6zKvQpnlfdDsiCs91s5tezTJyTycAg05qswSo9JUb
6aOz3H5kb3AxBhElRRak/ZXTjNWLI3hucPE/OZK1jCYk9oZ57YT2UthK/R/CfVeK
0Vjb/D9fmrWmW6rNO0ZxbZ+XA6ongvQxivVBaIa7dr1B5f9quVUM+3W1yrKrc/5b
zI4ggryEBBVTe+TFXRUPc0zCKJ0QKsXwm6f06i6Hb+79ipOeElNdp5wOIQlg2F1D
fl+RNCTPyY/+pSkHJwLhp08bDUlj0mk8RzPQk2ogd1aYs3bI8Ao6ExGrkZqa7lAr
qUR7UCI58ublxF0RGo3xFswB6HL8ma1sjna1YGdB+yGOE7fOFtXQxvrgiBltf0nX
YZwvFOWKgiKZyLSGcS+BO5IF4T3pLrdATXSlBnDPK1R7F2W5Jta5e80bgNnT/9Dj
J5GnRBsuk8ZVZxoL+mHDXP7dYWvPFj4NfD/ovtmE8xWF8hD/uAmY0/DwHwlI320V
qnZibmvynpjL07G8qBkxONFBcDN4d/AsYUxqWMypUDoQFJjk43GAPwxUYVUO1VFM
CCWUWmlesCNKC2LAQzqLpryZYygakcCVex52TKJEEmhxC24FzyY9iukcOHZK/Nwf
agOxJ+UMijWgpIA+0r2aZPK9LGAYijp7c5PSIhJdZ+0M4t7YJbpwtYDWZwFT0/Ik
s4htU919XhEK2nQx7oKoSsmIS9ClglWWHBjAG4JJY135PCOCm24Kva8fnmOxBANE
N0UCn/uR3Q1D8SVXGNfpuLs2g9XXk5hxcEI5xIwRsyIiEQfZBGbUISfHt2HyHIEq
c8AXardNhxLA/5zAA4I4fTI4yLZCeCBB3igD2qEnciqDg661lQxvXnV/0yaOi1ue
EKLoutmPKDvxiCHzOyacpDSWfeGc28uTNEHJYTAM3mCWgiOvdgSMCTmrJqJeLh9b
UXwSEFcxJ8x3lQqb99NRcca07TLRbgknlX9HzSSmDBNxVudf7QdnW/Ju83RVvSwh
hOSsztEXw7Kwq/nmSr6xJ1siyVQ5ZDry50+ImWtkJWeYS5mJ1mPdgb6KSqZpWLyZ
x9FQD++zpgX6pUPcO31UAwdRFdTAWXST8pHuMX8X3hdjSYtN7h/Hda9dau7qsC98
DZjSgPT79G1pENmvQ9h9JvnBJ2pDlFRSqWSfnFdmIjoNmA2sHN4hKsvFVE5aFLQ7
eUWfqcpQWO6hwKxhDqSnpJAJhXXRRYTMpbdUDCqsmhNZeXDYTH186b8Q6TcZqUY/
KhVp2/RBzRPcw9n4uitxbQiYvWHfkQpiwEm0PrnVYvb0rDQ59JUNx82pDuJwh094
99aY26OiKjD5v+4y0tJa+8ZwXLUILObXvERiFtZ73aYHi7PfU5pkyRgTht2WFKqO
LjMoV2w/Nosu6Z8nSlG0XKZIks0rKq31ckuMOxB7XtXhY4T1VTD3LfNIz9ZIMuIx
rQRiHla/+8W7W9cSqiA8ijS+jk1+lM4yS2nJUEBJWjBaAKcBIQC5v5rKQlAmXDK8
7xDXt8mpxZoHUnfVWPN2pPzIYuvWnbU9UYfdKAG3d8Xw8e7Si8KZ2tDedH9jYuTI
fwJ4XDDNzbRfFt7aRH5W4QGIS2uwiHghORqZG22FYIxqTxG2Vg+wtp2NQdqEg6pS
Ki8mIpRlb6fDsiycH4qw/NUn/l9aJb6AWc2g9TkTkIziwaWniXSUz+w6bJ3+1zBG
xghHj/jh95sMtSSxU+wPXsWzMYNNDJVdQJTUOTtMYyF3qiF4Z3MZ3+X4W5ReBntm
3M1B2VQH62wdF5X/jW2cSd2YLLjjkYGLeHHO53zfMoBkBMeK/6QM0StwRqdpDx3R
76sysPqg+kxYKwLM/xRQLSK+sqX+XqS3i/odU2fpQlNH2ZDNe13go5YDBlOnr3Z5
/XkAMf7HzSVIDdMo/HUGb/AzeyR0m8d7FYNSz/RlKgBGdej85fePPaMPDqhUxJxp
yMqBmhnKmldvUPSkKEvgUmgEOpdf9chAV7nEvjc6DI5gvo+GDPc2EbnrGjkgVr5l
BK9jUExWSNDZSMGX5OiY5Bii5cW51pNupLXLDEkIjcY/7YHRn4V1/O6hLC+mIgNQ
+xjBkda+cQV/pbbKxf8kuNTqimrUmWGehRNU+jeWBQDq0R5ueeF5huTe2wGu2NaZ
jxkso5ygXXyiXryNqnhYIyO9kDwtJfxFTkx2OTw1HMLyJo4758mn+pmvj9sUTvzB
SVsbZk1XYaz+aDZ8/qi5ntPNiRF7jZ2Gx+hwbuxv8frVf8EsVk9B+UD8zewGe4w2
KKV9jGWwdsMqtHX5zELNHWkLnYWV4vUOPeuQwSnbsbc3sr6gzw6w5/F9aLKmRklB
9Y9L20DjNYL/QWPXP2lMLPXGZOM6DCCxZSmAEZUlbnd3o9t2W1jIvQDSqg8lkEk4
gOZqagLjiQ9stixqCOEENXviC5mTXamRidYkrqOybUp7PA2MjdN3KDk6NIxcRuW3
hWW+69h/goXxXnHk00PHuat0xo3dQ83AaRO6KTTRdiTpD9Wc0OVJMVfeyQ1Ef3zJ
W1IKioUl5Tq2buyPeKzirhdXck5PKUySt6bAXjpYU/nu8Gaz0gT/291l7+Ienlor
DDzxbH66s5FgkKaLP02T8JwsgZHeraQiIvmkoWOYrpc7ko6P932VCGL095Sq6Y6Z
O506LSWsztJa0DM2mvlajiNuLDVyRD1oGuefZZEoLfo+lVkJL2hcTuxqNq0frnrH
ioFnzmRsuE3z0ARgjKXT1+HkKPBoyN1NaTOLIJLWcgiSpi/b4uiM5nTL5FeIUUGS
9YbZByu0sn7gpdNuvnM53VyVfzjSvslaZhtVokYZsbxrkpLtxxv/vW8K9fiKqV5m
d4+FwBaAP8xXlG6zSI21Jqoqnv64DolEzycM/Ki288w8fU1UiM5h+P0sN6nXc/+z
O1rSqWAjtayun7m5PWwz9MAtfi0maWiOuxKlAC0lTothBxi+oJUzp1szDjN+kVrQ
NP98+c/RZgtICYPg6F4mMM5eGvoSxcydkuSWfczC7vncStz2Wi6Fc/k+taDAUuZv
jZfCJnx+HukhHrh1QBByLi/4yYql+qg7KJ0nL7vu5xyRQZC9KSFmFO4A2hdFJj1z
iilsqYiMg5Z26MUKoCas5t8X3FfdQzKRCiXiU/EZH8N1uXoHJ66Jt+nuvEciH3R6
yUUCW+zHkvz07MStQ+oWWSh7vhbS5rQtWLIubGICigBl2XHuIIAFsZYyB9cMQgd0
awtVbJfcqu8uiwOGNshc17KIITMmViiux+1eBE3ZdI+YTY04PEw1L1DBl8PO7/Nc
g02Bt4M1jvYs2iHq0Q2iPJEQrHfM7Q1gMlIhNxDpt2A=
`pragma protect end_protected

`endif // `ifndef _VSL_REG_SV_


