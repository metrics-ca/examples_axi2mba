//----------------------------------------------------------------------
/**
 * @file vf_axi_mon_sb_cb.sv
 * @brief Defines VF AXI monitor scoreboard callback class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_MON_SB_CB_SV_
`define _VF_AXI_MON_SB_CB_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
FF0BYKHg4+DcF6GZibEfQJTqAeN5oKQ1TnnCLw3Wkbkvq/q5G6s2Eqo2G0qV71D8
MDvcpW7pZ9ZeC8XyEMuQxoartETeH2N8jSUJqZ2oKHlvBC4McK47IS1+jdLl9HrL
2ds2XNWldG+Y7Bkh0fXB36MLBcMOfZkK7mYbr6TemCqHwOQuq9cyamJxBuZ8PXQW
qNjM8GM+5wQpOJKKvc1VHD1t9eeleaegUs0P9fuwyZhJoBbR+FOhYo945IhPSBll
Psf1XOjY4Bf7RQVEXGhASyDvTSOtIxc5xJsaUTKXh6VRVx9W5UlimI663BiMXaWH
k33p6gvCAmGW6WbV+B41yg==
`pragma protect data_block
gqp7lANJQghnOb2iH1tR8XCpePU3WGSrcaiKV2ajxRIdPqNgAFxQPzu5chlum6D1
74K0rlnpz8LMP3042KBx1iWSt+WuZPuAC9fAP31IkihLDGlPTQjZ9asAXPpU5ful
BlNezYyFsgGkp8s9oJSaNP6HOla1q5Gbxu4OjKFsPnmUj2vQMPdEMZ5ZEfc/+Fyr
OaeOqcUeYnAKyLhPqu6F88BhmpIpXV2SiHHORDTp3syT6W64zIoU3hyoioiY5HYb
VFQV0ZU7pPzJUOOFbQG66HsoqMRAcdwxUikvizGr5pFoH0tVWud7MhayU0TyGM4y
hQOSWOkZROkw8skWqZeo0ziw41cLI4kZRILrci5y+S/7eLUssVpCk+Bb71jY9vs8
uNH3ox11YFNPWShBVIKVCjWWSv0waS7M+PNvapp28EdLNBGSyyazEMEqhP1r0AXh
D+qbCslzud/PknG5ZW7IFtHPNioL+3GdHqDcmG9Ue3jkti3x0CrFnstqc8rZ4leX
nWxSRrnA5QNoENhvqHt1hRpXUgm77mRrN6w8N3g9SDuiD7eUUQijkwinc++DLXHc
AaMY/qRyNLcUtW2A799yrQTVApzRtOuw2CbL8mgAP4M7A4iuGYnGqyhj9D1WL7Lz
OkotQojt2lezOAtwwaR8Ofws1S5SQ1e6IjUewblhvOHOAsYb7zJJcqESyPMg195a
cVfOCuXyVAJVYWC4YVsOjmONKzkKqJsoK5raPSzf/btYpTYF9gCm7zJepTeeHooj
S2/E8Ce8kP2mYDAflL0693V6INzcQKtr+x9tQqdFrsOsw/ElntxRphCbV24YlTEg
JECJi3BwAPGSjQFCw2q5p2YEqYZQX/e8IMAIUaRIHdPwizTYcNwN2gIcOMiHqDBf
4IUmImmvLXsOgIFTs5dd4mizemblQ7OUl98VeTH4NyxbLSr0DaJ7S+xYJP/TlGzV
eD1vuSftm6CUaJLwo6ek8VO0gN8AD4Bmo+OtV5CV29c/Myr1OVErmqu3Iw2QNkCw
rPX0Um4owbQWSfO2ZTNjSd6L4SlVrG9bHxjhCkj8VDMEOhyvaOJNkV/vQBRB34GC
RXAigHzLWvRibwd8IC+OI1Dyxs5u52Pr3iB7XI08r/amJkK0JS+ZzofAmhdm4ljt
IluWVXY8zZRZu6zbEjITVxNeHo7W9LjP64dcwv/hkH9WxWg2Mt2iKByB1dv9UFaX
Zyfivp+xGb6VlzbKoPD/L8HqACBZsoqX9teGVt7LB8AXdLyqpJgk84GExhKJe+3M
GZ7qcXE0ZwCn7R2pRzVMtSXlSeqeo87KSF3SpYh2pMk2pcrAopg79cVrH4k9JYf4
K+At6FfBSDkmWO7Cz9hcVg57oi14TyEteU+rLvndznYx1KxoTzM3Qq5YEd6rxWOo
gxH8d8Kt0po3M3sKAq8JIUqR352f2ZzaVM9aBa6alyVMQgNGtd9ePrbM8yiJdRTJ
XC9g0PmuyYtES9FDCgM8H7GLWGP0aPd6jc9y7wfFLe5Hg7rrl6Xct6MW1K2OvtIy
6odfdVR17v8YwOXuFjkF6uSyKh8Y3pRG502qgq+F86xp6tCCY4uE6VoD9QBvVcwz
OFKPCVecJXUB7d5jf1i7+UEhtxJQvIlrun/EmrrypBc9ETTjQF/eNzpSBtJRoULu
aQheNLKzS4Mfn1w4lcGt1zFGdgSqdGEbxWl0/TS0Ap4bTVqIUvIsHXzhpsAFAw1/
o1w+NqgWF40e5swqVTnjdUI3c30Omz4XuR8KZOzIcdap29/yM/XYrxAr0ahF8dMY
4lcrZkzA/sVWulgMv9E0JbpGbE+NvTQhJUDyKaLFnBT+Yy31K3FUEVTXD9Klx7rG
0cEI/gMfJGyv3x2bU9luV0gmfcv61SvbRr9CwcGnNr2w1t43BUzlcZV4Pk5R5lJH
3bp1/YteQzb6Di0Zq/9K3uVdehISuerzZWVyk7k8byL+Dv2ntC4KkdTE/MDjXIxe
/gQDuAUVqBXaKutuk5E5NbBxphz9/BpfNNC6WANpEh/4tdFO8egHmVodRvtJcGAs
lyEgGL0YmoqTZJTGR5WycSTzxO0345//53OJ4d+6VPqTE8tLquLyx65ts4hvW0E5
KBfgBClymOZDjCC4gca081gaqNWWtVMMGzx1XdJEHldw/1rm3UOh/l0XTuReNgn5
lhz9YYGnwXucTHZx5s494KvMfoUT3aDDeUFzQA4PrhwGjdVSrh8eQEsJk+H0lc66
WPPKsd3yQgozTWReLOpRM9Ojce8/Eo37Maxzuiiw1xBPvkviIxdnijKRO3xtn/tD
LQN4czz3M85F4VCQjNZe6MVwo6ciJKGs2Dsx0jhltvN61sL+VomvCNLPe0Gayv2s
yc75OLFncqiv30Bw/9nu9WvTknBHrrK6YeOBX5KxpKeDMNvaDokgQn18CkY2/YLS
HRnl/QwtKfJJuWThrFTTcPmivXEFNQWoRR9DUfOIpQbmL7D9vfEoH3iGk4UYyLRg
pexbKCYbfAhaM8wywsE79ku9EzIic4hBbhxq16xspwLuN0O50mHdl1RxITv1S15L
iEU73R+t8Xjm+GR98c/6mvDVagQc3wwwwMWl9I8azoaTOQcmDaVZ9q1Y80FFZMGW
lAimvcZOjf1Cafo2en0sGMaffrewBtArahvm6nzUyhQCEyRtrHYbhz3avAcULkgk
WtuLnv6TtNg0zVDgLdgEXeXZvZLGZI5ULQBZz3YkLvrHVs/avEBWLdoOEp+1D8V/
T6dQGBOoI4vjXQziSngpvwRpvnu9V/fHvVE+oFr8glKaNTFeZx5Gtt0LxtimNN62
6GFJHWjf9q5UPp9iRilXhRKvyBABBYcN6E7wPrZel9AXblMUZCATacCtwLwFbgR5
I7N9PCXlSUjDnS3wjjeDtwNwAEQEyxz/+dJhsFpy3woOdU2I1jyTLr6rTDpkGUWb
mRAyhKoRt1htSzt6uVezX8tLs52I7jmkcfFXqVWbeNEHP25hAPh8mkSNBCrg7hEz
EKI7z3nD1dZtNtTOBtUTaokKojQ3ELISZbBfh7TLcMn4CvNFGw8ls5C0vlq4WSlz
ujxVGLvE8j9g/Y+qQkbor89bdrJHsujEP0xFarnQxj6oGlHrL4owQkGh5p5VRFxI
j5XfNMwTqDfcZuLbC5GpFDl1Lw6f0rTBXOfQ1KFh7SSSy8mgWHEbUNMIBvUwxT1T
SlNvUAepQbnq/bCTI0Rip1eHiuxVZft5mOhILY4233zROeYUs6YIUh2ektqW7JcK
82/9LnyA7UXFAEFkP3dPewS9KPcFMF8QLEm22vs7UYC+qmo1NMwYohzs2vmGKJr7
5Jf6g+q2wJkDpOyJQQ9M10y1Ize/+jJ144kdm68SgIyAV8bCghA/tPgGazodVEau
V+OFBlzZHie1MbZPtURYLU4gJfeeAfkizyTJGZ/QZfPWL3ih807N6bynu0N890Sh
fgGjfeppkWRJkChUwE1fZztd/qDIRJPs+NVuu3p4qJaueq0MbcKuA4J9lZhp3tlC
lOy+KoCa4K2Vd5qN6qgtIjYDjeW3CwJauz8s236NTVaO/YyW80+DTw+zaLfrqg+x
eboaQqX2/ojj/lQpDZY5F3eRnRz5EZ38/ht8l5urHZ7Bug1nvGhx0iTQmPfW36wg
jTjDpY8VAI3abTGvOWwHdp95OwBPPLotE+zm9B0pOBNBz8d2UMjy2BguuhnLCqyK
1bQp7PoGFyauNFKQeGDeKVZSkFFsGGxVe87u6iWQgGxYgN0f/goKn3+tx/MgAkqV
7y+k6ECCK6YFD3RecOat8QLUdcP3TW75bkRTK3goARDUJUlV+QrgBKK3lo+Nx35r
MS6ziiYLRqQ3864ArR7VxCVyvyXGr4J3TRhJlyXLNHpIsdjb4Zovm+N/IKugwwod
iPtDY1m5jtH0WEQFxRjaID8qGyQlZnwv1aZ5sU1Tv5wFqSNtAG9lNGn9OH2eBQHa
faIS8AwO/Bt+wjViMfYPkC0KHhHhKsTCYk5kiOh/PcfweVykFpnbTooEHJsNFv7q
lOueDLxRvlZ2uaeBL3crk1u8N9sWoIGYPRIrIj8aLmeEysPHah8Ok4jxVcWkbdkL
75tlVxlc7tRiff88nlCjxs90T4xHR7TFUNNB07j0rIKs4pR5llNxgl4yQKF4UtQf
93ZnREpOXe8pM4KeaLJ3h2UjtAo9YJ5Dou9sZiDGFYpZWxaE0V0CSR52f1vZ9A5t
W/By/ousPd4dOPV1TkHdwBAO9Us50A2ygfUh1+K5CEwaF+gQ5WkNkuW6sXAyCK6D
1b4TNrf/7nUq6cLPUSdHzaY64e58b8DQe0dEVASVY5aFYYSqrN5s0z0tvrBF06ZW
qVJ2yqQST9Fx+Ah7hbNcrdpKrvB2N9AN8WuDfBGRCU5uBL3PjhUm2Ty18SORSvKV
FfbiklVYRKnFLUMgxkutFqGpqbWR+H7VsizbLI3ZGjhfpONuNznJmrOFuN64AsHm
KPzUZ6RZjmVLSfn5zv7AHYGkApGVlooPpZkyIWuBs4zFyrvD+LdDsEZOxntG/mpw
cpJzTqOQX4MWWfA0Au9i0vQlhi/Jc4Rc5jr/mdtDhsUBP/c8gO4YFq+oy9NPOefm
rwGuwshstiNLfKugRTOHsR7WpgIh1iK4Zbg15ozdwjXbn1nwFTlXERmtEk/GPpD6
6i8dm1qmjt6oueddmYk3g+HtBCF40JqZLV5qBmtI1TEmhJBUq7O3GOFFDgfGjSSb
iJ4j1x9xBK6l2Qy/21MVaqSBY//PMcS1/PkN829o+hfZyiUbyfGnsFXiXtpBHo/v
RoU4vsxv/1Fo6MgnAUcCOU8+Aiosv9U5lPs6pZVnvPFg7Lv8TZuqYDkygmo7GUDx
ofd1LZWxPAazVbSParUSRtkbbo7yGiyLkvEZ0p//n8Def+aTh9fbAerwjyYixWJO
+WKIA5q2UG2SChGJJUoIxAgVd8uD/QFm7jJkGrCHwVUqU/23awMsTOjZeouQKyYC
kZjKW/lR6hgMAfZPVtzlv7uS3hFfiRWkma8hB956NSQ/rcyhvKv94y/TCbkmfP1y
zxvqCwTF+jWeprQOSIwZABa0iH0LHM1Tvyu39h0gjm/CHboj1JK1LKXO0urclego
VraemGArYNsLj5oZUzq3ttLgevFm+fQdoCC2GN28DW8U8W+NuB+WMi+bcV39eFWM
ZXWyspuvLat9D8gD652iXbUuccwcLPM82/vxYKBUsFOLjUT/lEbfPJrO8Uevk0zH
DYcIW4zzllWYoTEJGh5tRztqmEItU1Ar7Y4HexXOwE2SJ7ZFbRhkeU/bxl5E3INo
v8UWj049UkljE39kbeJYv82mC6M01HZlFsMK5q7BU2c4UZjFETRTFw48yk3JYzIR
o5dAwBfMlIWYx3+PRsolgiXMASNk6vlmSev+87bXvNZYQWAWZKSdgOq6P/iyA04Y
V51Op3pZYZyVBuQWb2B9GkA5ZN3sBSzyJfxlMMaIawAkszXlYQFSJk395v2SI3z7
Cnj5g0Tty84rGmgZhOahPlfC/awQf/4FUWLZfka3TA/HvHt4okw8qxOiKQvoGnFO
HvRVZ0tWO+KQerlxRmHJduCCtyGxz+Mp9RP/sbYexdUE35ThnMfUrYKIUJEyXk15
ZDH9JkpRf4GIyVuoLyg0tDTSb9OxlzLsm8vOQvgPqNXoO+r8uWatBargGQ984hzy
itDHrUezI0HJ9IXXWGgVm1B+l5joIQjbUVxQMMOFjBz3kv3EekDaQLuDqDEZ6bVa
Rjz3oP43fD9LcaT2v3doToN7pSJWgspu2hYcA4kjcBGXEK7vOMovMimtlMpGOXpD
5UnbsIc+RczQ0YLcmVlgD+o+84b9YJKkVxnDhxBFU9Vz7ICacHxKFvYEXk3/6A+N
ZsRPVHK7BwGtJLeKRKjBhn60P84jNflSp+Du8LfaR96j2dNnJ53GcFXjpSWQaAoT
BpV83zGnH39ZyW7XGdBP0k5hRsqwd5gDJjQUPAoWOhTnnGmqBZ81zIhnIdTTA5TH
QqY6ZlBRKSBOjP3adVbTgrZipxAfjOrRg0ecSgsDw5uM8o1bTAUeFYp/k8rFCaHM
GecFQOVO4mvxJvuCET7u7yrS5+vTVPUk9hDZrAeQ5OhvSkvUN6PprpcHBBMTUx5J
VwsU9KHk3j4eFnYGMEfcYsxfcm0yqmqS2eJ+o5wmc+uFOrN4tmci0CWkdnixL2af
JIB+SEuNGaJ0L1E90vjNqB6hs52H9MghSKk94ur0USKqRWv9AawBD54Auy6NSZ4b
t7h+m8TdVZ1ZKzdpMTijUbRmpr40UwZGEhYKgt3aLnkrwhkGxSOGcRyurlTajgtl
zvI5D1tYkgvRF74k6Tpl8waMSc02TENjuX3QEDQrRrCTVZ2ty0O2kvTSBZjz/jeW
CP3kE3ZuMYYFmABeNlijXydoZuZxuORa1Wv5Pn7FKOHQYG+532zyN0zvY7XnMgVx
F2Fi4EX77Ebcr62Z4mPBDspKf+iTrfVPzBdLfQI+05Jsy2V1v/YPzRQ8nStEoQMz
gP819l4cn9DPUvNsAgV6HN8QRMzTZvYXTvGpBRCylrTSAGD8GBxPULv8EfoHLQ45
9zajbIEg4eVYDfWLTD37BvtZO3LVTvoo2/c0Gqobcpg8WA9XrJ054uyv0R1ZLNol
3/bUvrftbhaPuzrInICGsoUhD41+rMBA6SD8/0hJdCUsQUjdth5Tq0af/v5hOcwN
3aFtIEKhzXSB4KEErzV6YAZjt5Sn/4WgeTt+z4fptK1AeuY6boNASBNQQfl+UGZa
fQoqpsvHwAK3VLDbsHSQkb0pcRFCERTpg8gGmIZ/Aplq/NbbBByhmVxzLy443aeu
KPUnmxqwSpTkewM/VAz+GpSZgyl7cYcNHkD0u8aI0KzEO2AklFoIFghDhxNcTTqi
/Xu9JKVRYC/WP0JoMBo7n869DKg0Hf7khkdFXoSuzxrTqBi511TKegx+bpdMUl1Z
6qSZaJdKznRSPMzaZ3cP9huIo7Mmifc8Ami/hZPWHo+FSQRwpA2qwhSXn/I953e3
5NFgLAcpozHWZRUNuyCkDFqREpKFSdNPP1+zqrSfGY7U9nPucRmDLGq/jKue+Fde
tByB8aoMS6kngaIN3sVkKM/rxuTN84dA83pB6ty98bni2IIjM5GoTWt/+ov8p4xd
d7n83pP7RsjZOnecTZihX2MMGwO8xMWto5UNZQIZSIH7SKsVebLBbPh+Je5Q9oek
thO84f7viyF65s0mjtEiOlxQKe0QuVqVNgJUkbi+gLw6h3UVYlRj0UhH8gSc29iU
b1ZrNzK9DsZK4q/iSYm4MxM0hdDM1U6tWGJrgDXQEMwAidmFHk8qo1bKZtUMnzHT
Eb+Yyuxe0Te18zEnhpgKfQ1V20jqx5J3XmxMZAowl5HS27qpYKtgaCNrhreU27bH
hakqmqx3Gij3KtOpPJ+q1QHY2DrdYckGceD/5iOD7sV7RfK1ucvfWYWMkDmmi0p7
04dYw+R6x76HQ0Crf3BD/zC1HXfWIfYk2D6W5db+fxQnFNDTq55Ac78j7xzivUeF
i2vHYWal4rOmMo0Mh9t4RaXwGZnsZLU7djiJRCHUoZYsapb7JCPUFkspupvhPnQO
/lxolJggEMcobbE71mOzx6h/kQylf7bQywu5kfv1EwhffRc9aE5XUHU8vLU51QBN
gMW0kGuwZLrFEnMKDw6qzuKwAKgVAVjMIhQbIHQt4+Pl8eqa90bepKLrGPc0LKld
xFm6FAr28Whus64sdvL04zZCDLHaDFNdsr3gxzYuk8USR2I+g1yeNHQfu3aqCSaJ
qmxr3RW4gCo4svkKYKIjzxtll/Fxwc6bDLBflfYQqQLMyQ43K52U56tRujNZ8x5s
PcSSfCtTXD1WDM1IIOfbt9HjX3kXbjFtKBn3KkLhx7o9ep+N4MbHj/hTqdG2ni+u
RQyvyYe1eCCZZfJvkzAbF6k5oNhJB+TdudRXo8emK7TAehha2jo5NTf5MkvUA/R5
gOAEz4w3iW9+MHWHQw//efVsBNzv/poyB/nioh2S/YYHQEclr0LifxS6wUYBcW7J
vHajUwvGbqKi4j1g6UeJ85Ce/KBlPxGVZu4q7Ew7QAzuEENdC53adMn9GoBnlY+E
nk3IZm4Anesp/ritTnTfGoqc6Mnm0OO/HZlGrZVdAtPekSI7cuFBc8dCZpf1Wsi+
sllf/IL3EkkjWyRlxG6nNcLcQ4bVrDitcE4QJbpyB3g8jmTohGW4RDnnZICOd3x4
4AzMkiz/PTSrFdkGFp212W5o3fHmp2y6wGmzOon5oK45Nq4E+hRKfy/MXeut6toF
DsarqskrK2LKB5DAdCWOdDq720YAH4hQRYc7UWcdnktwey6FgHL3n2cnbJBxRTf5
S+jKNlgn2xak/Nw1P42vF+5J+rltCowArCqUkkbCekICnYGaTMfmT3knnegHPjAJ
yjZXoNUa4f7nlFLuNAriSbRgBJ3DN6/i0emljBIFbC+66KqRA4cNq3HNCHKvbrzv
Rh5z6bvBiH411y0l0oKlaZVG2YwWUnBJouBZ1x8sSoYC7NpMgS+SXp1cU0pLGJRh
hzwq7MIiqESAOdGfLV40PY0zApd3yv5OnM1PVEDmx++q1zyqJtlmZtQnX9rMrmZv
hruvFwlTGFSqQFsP5EUfgsJv5aEuwH4vZY2E19zdkC7rXVvXRZjqcBFf7o5ByWtE
yKJLdb096rCxqKQPO3qTR6GeH7RzjqWXPv0KCl5PV4EesujpFOoFZlpJzhjaBoW2
RV+7CYCPKcWIhnBX/cpBBDygA5KiZqRLyv2mGrGhOwHF0Q9hz1wWuLnmAuLRg35X
UYCGp6J0G7OWBC8y+j6nq/GrUAUte9ir8z1wjm10TwRCd+02hB0x1kMD/q/rG078
Ld8v9AJTm6SNifNNNCD2ZxOpWWhyWOe+bG76ZGdPBObcvc7XYUCsFOt0bj2RvZkH
7M9AVBhcxM7k3j8+USVwEjqmHUGur6ySzVx9uhd7zOpTNupHgwMPjjIna5v0RWSY
b2MfiNDJsGO9mM4b1tDeVnrDMyqF/Ui/y1wWZSkXYjpW4bxCTN1sQ53UKSoHx6Dk
V4oT1NK+98HIxBw9hsIrG7egmpYsqdhPr7u18uEvtHxI4sDLC1/TNuJkfHAemJVq
EwP8uFs54wLX93krTdlYv9Q8fQhc2Rcqy2v7ilt50fgsXaPlobJLQ57AQjfYnDmn
eW3Ltx1yukh0dOTgLVj+suAEzjm+tgUuOcmCJCa0ZTAeZTQ+1ffWckE9c8WhIZff
Su8d6y3EmCQpQA3EQqo0unYAGqJobj6ulWOpq1cbuTDeAMqbYDootcP3xrCJNn6n
wlyPNFALaIe7uDNp9yyCQLneWUtkUcIis5d2gIAXMQkZKkxUEegqyZEAiQxtRSAq
kA0zZX9dpAqlXiZ0FiYyCbGLCwbBcsP1aUShKwbx1iOOZw46FkeBYjoIzv8WPEfM
H7ujiSgiJyD6NnyESQK4uYnY+0xLvBSyjEQVTtFkVjUWdWlptXUPV5jdBAQlTKDw
mdsQqDvE00J1tTFr9AO3HYRuxZb3OwSzhEM1H8Y2zbnfQW/oHem9nPy63zb5Z8IC
Rg7ZyvPqH0eK0FnpJKtkQDxJj1YMJMHzEcZR5RGAwXA0rQPSlhqnv38MEzQb+GO3
xKzSBZ9zM40SAbtqlXrm0UF09A6JOME8yPrmOBiTfhRqS8OghtAFIrtrIZBk4hoe
XMlMpUsynAkkvXNVlxbVoH7J0xrZTxHEemsxqflMVmCgGwqKYyXp1cQoYQW2mMkx
PaKq5usB+KO2GIu9IoniJITpkDfBP9X3cbNnr8iwOIpQ8IAgnguUXvY1lCEwuaAt
o8a1bhD74t6X1Yk6/ZzOgjNUq8J5Xjzc5+6fRpRa3ztybcfOY2FmCCKZiw1p/1pM
zpcAO3PckD9ssATIgb8TvDD4cDQN3zg8ESkOcGBtIQgvFNy6l/M0jSf/iRsHi8EI
2oii5gFf4BGVpplQ1oc+ph3Zb0J0FaHDGhUK9OYYiMfgh3j6Z94JzIAvTEVuBimb
w72orWtyAkyBaQrtR/VqjzngAFo/bRYya05zlM79Dqkhfsjjri2Bm069Qu2w1WaY
zuPZv1LIwWegFZJ+jF/KbIamfWJ3IUT0s/AOhoy+0swxjxkv0utF1XwjJBqF7Rb7
vAHBb7V51iMqxgMmjNCaOpYRIJp08NpSUnzARWuEUBUXqTUrqlUFo7Q5mFb//wHZ
`pragma protect end_protected

`endif // `ifndef _VF_AXI_MON_SB_CB_SV_


