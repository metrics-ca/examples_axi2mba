//----------------------------------------------------------------------
/**
 * @file vpr_mem_typed.sv
 * @brief Defines VPR Memory typed class.
 */
/*
 * Copyright (C) 2010-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VPR_MEM_TYPED_SV_
`define _VPR_MEM_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
DcnhRABWdRrT/AdGqmLcOPuztU/qMLWaR5SGeCwRF4xUW4TuXadCGLxG6pCgQDqx
vWWceo6LVCY2lBYlzwSTOfLe2LE2xtkhJIXFu4mo/rjPLZkmS+ZO4OHCIQvqhc4R
Il6/qMQIDg608LwM3HIe97O41mIiRBmQwjqKb9SOtFCCHZMwVx/jvtOEPSd7YQHv
vYG+bSikDIa8TG3rxBI9+9mKXhyCWAM0MAw9jK9pi24N6HtbA5b4XEnMWalOqWZS
VohOh0CkTN26UNm2D88tX+zAXITk7HSYgUXtDAOTt5jpyTeiuN4OdjniGGrs4P2X
4mLP9wbLEVw10mRbdjSgtQ==
`pragma protect data_block
l8XZbEbpWb9stfdR2ZR4e57YYwT3ebyhAoMtJCq07BJZ4IcIqjFPIaxirqoQ1qR/
Lp3qBe407UKC04fMc/4JrTQTOqzLAUzhP0IdKFNZNuXbkWH0OrDyxodxz8zntXlS
DdOYTek1rstzT9Lvxv7eaEwhSuuGr79KMo5xLV6viRXM/2ORfPVZiOu58ute0elI
b/GvO1sYnD2o5SikMmxmh+mlbeRdbgReGqHUjyVClj+lwNADLZIIieXOxl5t2Ayh
GADXKn/ZbTEcp+jhp1W2UGl1ocBzX2UVs/MIkiUoeaTaV9S6zIEokI/y9iK3D0wm
Lj2k7m9uqE6bSHAnM1NPfMXZxoy6w92P8p/2XS0Ef5ScMbe9ppAq+mZ5rgCsIKWa
8BPHkzX6yPDQFJ8ujUkJWE0ISm2tae8Jrp7lzbO/b3/hGe5DTZqrnsxfDt0gUPnZ
Bq1uLIrjrtlmjj0IDkE5Wbh/DJEOnMa0uzzygTNthZvNAlPeAiIWxFHYpvdWCKYb
DMSz63AHMdf8Zl7DpHE8OC7BT0SpR/EktUpsncuHyPmt4PBO7FxxK0bnRRMAgv+5
Tr3ksrONufCA12XzIzHVw0iH2l12eWCKDVDf07gf8FYS4DkUwzVVEOUGnGwgKCrI
WLMRAAcfWm2eIyKSYgb+BooK6R3RhsMWWS9ywhrfNytkJIcufNdw1SRlQRNQRG5/
mt6ugXFpP2ZHbWylnY/34jKUeztUODf2HfMRtUmSr7FqHe3rNTfEvFqI3KMM7G2N
k05RZC+ukx5axOY35mGmBA/hWBkUcjsAumBNuIBPGRs+LAwiYvaZdHm+Sc8jERHu
BjJt/+xt3bqGx0QBYZHql76ZKW+LWgMebmtI5heTaybcMeEIYx4o8I3RHMmhIw6w
lnOq1/IOoQ7wd+ljhnBSce2ZR5hKoJlI5vFBy7h/Xvn5g/IxzK6tvH9E7P8GEMWH
NlMFpQv4Pvk/2JQdEvvQVWNn8ud9jOBmz2UN1ELTx6EDI1CkJKdohxQfkKrsroBx
MpTHleqBqhCY63GF90rZd+G6LH7aNZJU4GtZFGVmJySRnqmtsOGcA8c2t89oKnBr
PVT3kkjxE8M0zSQpYekAqyrZNnLFQ6OxEhoId3uEN4aATC0XL9GiY9tC+ZC0NF42
ECR7+WTuLkiL3KYbEcB6ug8O+r04/v6H2pIMLmIM2MO/D47khGlHODVd+ERDAzhG
p7UmxLGzsY+DvlYN0dAEuKc55qpV0C/Ab+SgNaLVCpRx/s8T5wDVF4wVvb1WhfuM
C9Q1LUTSZTfCk/GqIIxdKYtXI8mkPrtpgdo+MY0JSbz4iy/bamRGI+4kzyw/nQPF
UNUsIcF+77oFP2Sm1FQKJjWUMSe6VkytcXg+XcHqPNwRV+bh+uNnWBHIFRJ3HZgK
kT+Gp5pYMV6+vbZoL95gutLxtXrxPnYeYMM2Sumrgud15aPVBSA5POf8oztgXDb1
3zVyRQLa/BlL53vFC200wezw4lxyn7vSbDCk9J6bAKvLCu8N4Minv8CD/wxuFYLp
hPhqTI1OwvpJuwcfEENAic+npQ/wY9QY3TRiILUXhdIexjIIIYKLcsPs6ViMP4OQ
k/IRIkqaF2FToxGG3sVLsv2vY8VnZS2IM7qWHWda7Cm//oDgVOfnShJucI4uij3L
7+cBXKIPK2AnNOhNlIgvc19KLsH4e+UXBk5P2Tf27C9b+XDnSbk3a20TZkUiOA7Y
e88Ggj8tEsJnPbVz3El8cdv+RqA4NMIq+Wh9RspYRs0wZ3LSUsUayTURb2o7vHFy
afrkqT+zS8O5V02DX/9lC+Q/mKoTvuSEvgF7iwAom2WkHY4q5mFLs7zPQhPNfDW3
pqBUTea93NvxQ1Dvc15lt6ANx3O2DDnj1WVqcbhzYnC61HaTzR4khVCT8HR4MgtL
CXEvjx0VHwsr+R6Nb2NZwrkwneLkyi2wsyDzSAhdEToy+7bHqbK8UGawDImziV3E
HGC7IzUtmbOSbjREMI49x63WeFP4S0pUVCT/3VZLt4C86D4N6Izj9zJHC45MefKR
zY9ViQPr7r8DtX88aw8MYXMCqyrgtplW6AiEUm8Gh/Owwqg+3G16+RuRdJVxiaGi
6yO2sVRFkXZxdpLWns0Bq3fw08kr2VZet+pvIthaYKiPK8uE5aK/uGmib5UHoaT1
B8qrVKWyPa1iJN9jtdq4+LFXQSe1/iDFCGugb4m6IirHhsPpIt0HecyJAfdp0he5
27bRpF1c/ZPlHCYXWNZqYdr7/OR07C4kkX5+cOEc3WT25eFP6IEvc05Lz3qHQMin
pr7vIxdFZwaOfn0aRfPuxCCfFPdwXQ3/mY68DBCRkfqiok/wUXy6Ch/+3YMbaLBZ
iGej6N9YmbpPdrxTnr93kNE1oK8HDNR9xjldXEGZRPim3ck7grkRI5J3FPmFnxE7
RB6CxVhQQwnW58QP8juD2Ab80A14K4l2Bf+70sU01kKTUQBHvcizgDPQ9vnMaw9E
O0tvB6jbA64BU490HJnLPmgQ7Ce2qEWRWP02sHiQ56QVzOEL2r0+z0e5pK2XmzRd
FH0WzFfT/mM0r96G+oG1mXa4xAHuqHlW+ny6UmxEudbP6094EDeC2Q7baJw5clPh
ma0q0SFgeSAD+mRVYBEs/GWAjysdPDn7SioHg8o5E3gWeqJ4igmbE//kS+XPc20u
a9V3O4Et5mtUcRda4aaSIeBP0Gtg/U7NmtwW2uG4me+uKYo3MwqfhY+l4Hekg84y
0+aU6KlqFzicFDvEHTs61RaNEDzIivQ06Y9rY4JNJfVhtsaitp1V0CD4JdPIgDNB
Sn9sTgmXwYkjhd024tGxuVRBOKwibHaNd7WNoV6I4YHBjLiIIC3o6S/HFQnquM13
G1/KRUoScMRm9dNIWWiyzneyurPjEIZQFCQi2/TBq09qWY3YVkBjTmZ7hM8fMpiV
Mac95N98UN5ezbmnm0Mk8l6ORmbEf/lXRP9ppt0Z0n2yVeqB/b3UAyw9/oBwGZMa
B1KDpOm+OE3w1SBvS005eA7+EZOZuBq/3LZ/LTafHjdW/6SCHrdUUgfj7uC7UTn7
qhqV+zklXVAv5WpE9aid5LFmhRoZrVtakbzeuirfqHRIQY3SXGgj3h8rMoBfu92f
XuSmCuXyAiBXfq92FKq+owMKkA7tuW769idg421NesvbKplb72PcB7pA+RgyZT5K
GDlXwe1u9SKYUB6bdxrQVm3xCuCLmqOZcfsiMtc160EU97Laxc1PV45ZewiLtUu8
7BssSTaz/t/HPTib6dcwDZm3TbBPDO0Pmzf1LLfas2W2iksDvE1UEm3EHq9fOZ6a
w0Nowl91q8PUrgVMEPB7sOySbag/VpP5dWR8+/0wXzVjr7E4kgXsvEu3oM6zDUUo
rQ2eD/AcBA3ClsIYz14q7uop1QVNfj3JuX1Q2W1ddCf1NdZuRTyb3qxtq/Jfnoh2
BEVSZIC7DxBMZWdM12O5zjgUaIfAYySkDD0W/Fm8qePRHi8Mcv6blUQiysMHpXlE
pkekmlX0gDsmKhm2DWJ98xVVUs9HYSuiwlvtSbEPszJXVY1+3DV+HJJkPaZ4Px0u
oHr3x91c9Zi+IXMkrgB4QfS+IJ0UlUxn0xlJZMPrUbkkcAZUaRPyAi1deD9DLhXi
RMjc3AwHiQW9/10yMYwcinsM7T/dGSe95NOWXohoko7M1u5eJMtpr/w5b1VW0YEu
tT7nXenC1QdX0pehttjqf0edcisYZjd3fcHn+1agVWsqg3u/hLrlZKpnh5vsWhhR
D1xcifkJ2SqCMxklb6Eoo03yRDyWxYUaLXs7iLO2J8JtxvglX3dUtLSimQixhVn3
4zjVTPlZ5jehEI1HM3L5BffEu8VrNx6SVTStBZ6PM+BnLT7nJRwB+JPpWUZ7RIPi
/GHlRtJhL1udBBafocqbzScSdN+9pw3fKSILhAvmwZR+NGfyakNs6WubVXdlxpYq
W7/y8WfhgePEr+GDjd+oH+/Z1crD4nUWHHEEuFiCdgteMa6FOMY6F8aoJVhWtidp
C9f5EoO/jb+H7YelxyDLDLndlkIhR3RArWEvJmKgBC8edECv6I1yTGBXDRbFg36z
dPYT6cfsZ08BJml6RjsTe1iZUfJ1FwkAwjzR33OpV1aX3XLkDzvZOMcv3bNGswmf
elPRom7po+qCqGLIL1hFtcY60vKeGK+gMyPVnM6R0K4XVoR1htCkLCOnZ/SRhhhO
Iy62ruOBfbYhhmvjnKR8aAPFu4f2sGEGpPqWSDvFzreFuC9gypGGFOXqHhzA+gSf
H11WDsaenikRGf+w6qEloDXiTWEW60yaidKlf2CuR9Tdi2oSuVj8xkzYGZms0ZeV
Kq7bb1ozunSUC5pQFTo5uX5yEYcWDr4oIAQVPJ+XLPSBQ8yHJCSK+G1mT3yAbWo6
BiXBjo/ktjHZJn1gQi+nUd0AihpLHIN7VNHC0ddnwyWNI2qkrS17Rs6BQwMZQi0t
yyErYz+gX/gsNF3RuGYeRqExq+ZVXm5/uwtQ4rE5GDasyMTPMiqyiZDSm20I9DT2
GJ2GFqJpF2Gjl+tHy8YZF6kz3o+8WSuFKsEP/BwkwZQYYFI70aRSk3s5wk1MBo7/
xnyNVroprZe0mk9OOdbrlqhOpnz2eNdb+JxF/1413Rw+quSvPEDeOgQMfejFyKQB
60SY5auYt+gktPSD5vZt0Yh7twYjwU18gL8n7sYSzXFdbL/IdRPstz1PKg1GErXS
15N03AEyX5yVakXUEHmS7/0zudL1BdjukUsU3RVydu1EzxQuy8/JFvkFe2ue8dIp
XODXsFaDl4NsXEAycY/cRw4rm3Us60topbcVk2bK6RgoFD02XtnSlBcZoKMl9awo
86M4UBCbPhqZ1GX4zHBvVMKrugH/YxlLr4eN7cVLDRXc5aEQT0K0YmkvfdLrndJq
I2VLoZbbW3NbkXW/RjIhMD2Yi2oq/4i6MUd5kj3GlSYat/03Cb8LJt89oeX62H66
4unBU70WmwkPtYZcuavay1cdS0yiCHv9e9lOS1NRP3GTy+hxY+qLURTdaJj1B+rY
XUigbC3DU43J1bmm2UpnS4zCLEp5pW0RPixOpms2AJXVGqjHDiPIc6umJR0BawTf
qbRAj/vXG4+9dJEUfft5uyRjb/Ue4KC39XegZhRgGNZeLCdlTZ3CXozBp1AQsYED
uNiLXQNciMwS8aWwGRKTOpCC9DPuq2VfRAv+P9EJpkWl9mQqubnfkL+4/z76fPMJ
hRFZPz8pE5T+kFBRX1syWVRGOwiznCWLT5iWXzibfzngEs3AkmXRgQRbn1DpsoFl
Jfn/GBXJmsnCYK1TOPPo7gdPPRBjSy3xbe7QcrVuGDavjGr3o1yqPJ6iUXs/4dAB
KOI7JMcqvMqpcRCBso+ozJYwu0osworw0bkdNRL3jJhKshJdN1CwnRocXMbzUTOl
VqzDom3wxgHpIyFf2rR5iXI+btWeDuK9b7edw/JOcDEDjJZv+3Xo5H398/9zw2ip
ICqlbsEihIKLjJCQm95bkWO6rTcO3WnfzIaXX4FgHLkqp5wI6xKZVL20c5FcOxf3
Dfk26plOjbB9QaxUnzefNbgP/iNANkla3/L6yAY8ZoWiQZu9TFo/8lYDuSj6ZxgO
1+RHspjjnfcBUkgOLzJJ8QpPh1X89Yqvue/1vRHuOcVrCHdm6yHsTD0ShIylLBed
0tfN2UmKfPFc6tuDbGhgSky3G/WJAQDbAyAAwr4JGH8f2r8Ky13eAfFTTMYbBGDc
QA+6o9aN1iRjGMQwYrlfxF6ACABVVweYYDG1h+FLvn8hJjtOkc8R+lQgsbcBjHEY
gbq5ySfTGjgStu9SQVlDMOnx9w6Wu6MaJLNK3S7sdGWlICwVeCrpCaKNTDIZgmf0
jlkQdfGPIaxoiMds6KIMo40Jk0ApXAprqJfvUUzHIsita34rMpQYfjIkyVJTOd1y
OmmeeDrHDNhFVJByOfxClBaNUJNu/penQ+Nh/t3oOBEGfpXADfaqKKXCrvnr0Oc5
dzMe4YJlglpo069gKJSbTHmFqyW/yOGOchvm3ohSVd/PlaRqrSijbTjL4Hcl0hej
Q5zjByh0BBD4N98pOODeMHPp5PBzy+qbLWbidhF30TPQzHRO19G1eC3smmr9GA8I
Mbb13DJT0u7I+KTMsv/IC58gJt3xOYatuKyG4KYEvmIONbM6MwSoBauXoAkvTybh
xgNXvwQXZ3dSjIaugsKCLqeqBoHgIAXCk9MRUo0LETdzZnKJy0jrIPWy9fpmUlU+
+aCoD0quayJYfhOhHc25ibif+R2ww6pEhawpw0vRW4C+m4gtyvT42+wAw/Ea4bmO
X446ziV7Q82VecCpsdiBswveWUBVYfwVWUbNfsNYYP+MT+3fzwt5MaMBnDJXTbY8
5x17XDT6ZXEVV+wdcTMl38JwSxAZ4VwGSUdmUPia61PtUlutklMZVOtmVuhCFKYz
VBsYPoxEpSRBYErqiJx9s/TIkDaUi4pjPHpx6bqY+hWojsoh6HkicLpKT45ZNMO+
rVWz7ya1lK5ER+2w8s+KCacr0kcJuAHseVgYLIDR4YnyVVS0M3x8XR2Q3HCFtJ3R
5lMNoV3WgkqCtc5+D7fmWxC+0SDS/PqJhnwjNwlnTsI6i/btUZCHFOmigXJP6c3X
P6zjM9+OSiBShVgWIm3ISIxGFJEX3lILb8uZqkvnkFhhhUbTP1g0TyNh0AXjeiGb
ic9CI4SjTWsntCX2P5SUrGynMG/luinJujLcnXJnQpzOdXIHO0vSocpn/D6V7yQ7
mO5jf55gmvS7Gi0i85Q4KUVZjHruVUbO5W7wLY77w+UVuSatgj3SQ8wha7KBaWoU
hSGtRZz5y0K/vBl7BBdlNM6yONyfgou5MXrRXQ4A3Qol6A8TUDsQ9ZPHGGHyQvk0
hKHQm+eraEzaCBTx6u/rZSeHcF+KPtDDWjNp3+QWcMVztaw7RYxWMYkzzMdB+1UG
h6wN4WwQ2fW5coHTwl/K/XGN+cmoAkR9OSjjNen+odP3Lv3i2LFHFoVcivYapjjP
07ueVOLy91IXNPR0IKXq0MrdO34+D8TUI3Aa2a4ARBuq+Ij0jK9vnFLoSacRuBRn
NpbZHP7ggiJe9J99QqUSOc3dYli0FztsRsA5Z0Th/dKUvr2W5spMZjoOJVtzgQn8
ycEO3bee6PKUsSA8MALY+uS6+eYBO20YadqlYF4dwQa1anDZ84fSyqcLc16qlZVE
U7NnprFurwZfx7HEq1bVTsHvrEOOAK6LJ4mUbyTTnRY2fFCs9DtWp6wbUUyZ+cVW
r+oo70lD+dAiz0u9fhslad7oAk/gfSkDlZJUmHzdildL8Kj1nkKd6/HMmtDXTbp8
TWgAq8KsYGSgl1y3rUEyyUCHbGZS8BB1yiAhbUfK7OjTL+QBC1f+Jv6GxeyRLi3d
zQvn6G5xgwqjA9KhI9SNkDjbn4Px/QrDrRrLbjUYOvQz1aWm4E7vawQaR58tixTT
a7VN9F87VwvmBGDb6iccwV55OZuTdKKXGUK+a0Q+MHHZBF7zDAaqwypYSXVe6qRI
JuIVfkeSEgx4h8fVmigwJcRBs+c4w/QRnpE2R1DFgHsBkHQXs+Za6fM2kfRMel9Z
HasADZoHy/YofxjmGGCisoNaxdD5vVylZ+ekGYfChkSCbiVgdoMLN2mhm6rUuX1u
5gydieg/JQsWSrDD/BrOafUYLW9zwHfPQDSfTCXuuCq4c2rwFcvqsnpdyj+TbazT
k6QKkF7WJxlZWDmNDND5voHjeDY/Xqa9L/KS3QnTE15EM4jLxNUF0AqhrYV6yxYV
HFsRRoRoXtrvxL+8hHBpJPIUmUq5Pf8W2lSS7wA9dziKhCwRdGecrlEOQ1f3o40M
MizZgafsBbXMU780yTHOpQ0wjRuS8TTuuGknK30lBFyFHXdiDhrn/BQ9Olu8Nux2
roIWkcl23xaK6qkAGECF5m+fBsZuOSi8QHnzZCwYWrYBMWaEuzERhgIMb4yj5daf
mtCgkmXKF1Z8jcVu+w2SAEEgwBx48J3ppvWlqOFQvYp8FBlkt9HR4wv7jJcGpH9O
5xGmGxo6hD4biMn8lOJPsFbNBZcQQn0q+7AMXrwE0/wLjt7uGDB/NZ2OgCivyGoL
ktc6LWjgb1NjFk5JYhB9BrSU/s8i/TSvaAHp0HmHI/X2+nxHLZEkzqhDNI4UetJP
HcYeWZblCGsSM2vDpVjSD3s4YvIe5cy0UG5bNfcH+JmQN6ceE7dr0vY1pWamJMR/
QA9r/jmvXk6YJ99tnFeSCe1MZ6MQkhKLkc8Yy7Q/qDFcRVxRvsVctUWk4J17OEFD
CAxnfetnOMt2q7iKM7ujnTL6XTSpjNGbmksqE+u1S5Wai0KIF2ZL3TZ5YwH82ciz
zjz+dLGyNhAOBssYq8j/ThLzSLcmDWH1p3PW90J7cISbLTagEy30jrRw4BajWCCD
xWh8cQqLZ3hVOhSv17eN2TY4LVtBcvTOJkEukyMQeCcSaTklqjD87aRdodQu+kxk
pblABENSXqxYIoeKV/54BMy23Re5UvV3DF9kQozSWo7J5Y9XvyF3Stt2FQMLYFH2
sk0PEN5p18m+9D+ni9YMHNqQL/bvrObiI/dAPEEk14zryYyHgNjoLuTeGqcaTbMS
f2NdqSlGyWyrc0R2e7eImOye9YPwwxThxRueszqejHOLwyDJt6Zd45sK10bngaP+
D8uzXYHPghMRR72CXyWas9DfAS7Ri8FQdkTC+IpvJt4TG0nxpECKMuKbx8VXKSe4
xZ2yyWoyGn517oE1IfB9H0fOJ4wA0nHHL/rMTYgngjfAOI+3aeQCIqWP6FCkZESb
aaa/uRk8Te8bB/xcQ+e3Xo3aW9kKh5ucsw8NCsVHuctFvPzKQ+DhxpV3UTKyRuTl
fDKklB7HkBGRL72nIu6jQ78hH7tBwLz/ULsv/qmyYotMcYq+uTqqk3jsQFzqZExI
OlyOoqmzmiRgpYkJ9+vuFpW/8oaBed+UcLuxKAbr2rxtDVwHcZEMkZiHZvwvpuh3
Bvjm0vmFJiqYjt3CRreDYFzctu4b3eCmlhpI5c2T6mFKGnB+jsp6U/YA/6GpjsNs
NZXS3rGuSq9VAxbDw8LZtXDUxu32jwhePB44fZSo4Dt/HU96lKD5w32YNAIeOrJL
mp7W/4rxLnOYawJRpcHuH/jZ9i4D63FA1P28NL14FDQ8BRwazfFH+/FdZeTkrlhc
jxviSmmOBXaVENuBTVr71YzJ2R8DAqBgLtmPJ1YyEWw5TDgquBMPH4fcxNiUSf15
qMTIfUgzA/elabKbJspHnEuTDqJX6iNIKjf2THBsb0CrwQrTexyAsbrTgMmK0Ntc
gMYXlj7sJ//PBOJ4pEpM3m0HyGn7Qm7R6vmaN5EqqJknhPPs0aXvnrgw5zKefAPV
P9djXJG9s+Q2OJO7bzNXLO6cMFsjtsXAv6LHcVxBX24pcUK0pF0j3zIG8ZzDckZ5
blQVWBwK1JwlOalxr41oW3OB38ZiahqXSaA4xMlJqVswpYJWqfNLcwrEni4zkV35
hQkxW7cOJSXXI4+VbMsPFCHKeC1nPtr2L9jb278rNw404aod5WTd/cy9qJsFa+CE
Cs+u9QkmEoVmlmy3hLwkhyVyXedCO99coYeFkvSKAAx5WTJO4hDE3XNcUC89Iium
l7CS5we/9thxbb0KnnxZ1Raw0Vkyqo/Sfr3b4NcdskIXkVYba+G2K9h1rTAIn1cZ
wQFGsaBAdrjxqoUpWMRQNJHUiNqq4vYaauxqOb4ToF6QlPoM9sn0yEJEDKzKoW6K
1nSV10059nAkuR64Ot6w+wbA1XFR3yTq9POZaWEiLr6JRj74X2LtTuvlYMlBXmoC
5NJpoZCQJzsunahRngjaQ7FBuGv7Tu/Odd/at7ea436+P+N8Yy+Q4JS9Qsr2aUYp
hrqSuY1I8FNgY376fSn7HpGlCiyR3hft0vGsyMxmvUnN2TxGs190s3u3nXYZd2nm
0xqvZoHgGRAJUVEdxUcLkUR9WRlWVWOnUsHswu2Ke/uMiVF9biyLVDCc7R+eOJbl
OW60droQjCh29rz9iABx+0qCmDpIRrzlmF7AlSVQpWxNDO2VZghO1R6BUxlypHsY
dNAcFbliMuyB9MnDjhD8praGINksfVbEQXEEgeBLvfb+H++YYlrXmXw0rOC/peZ/
F+Aet7mZIhIt7i95rM2pXdw5UWUj9s/bJidZqAtLiN+TmRdRHGW7qnp460d3ZMQE
avgfithlSmAiaVUPnkd7r9P/W45+sxU3RYkop21gamogCDY6M2Y4vj7UDUr44FzY
aealHZS3C7rWy7KlzSHRJBwH9FbbwHbQe/s5T57DqJjSPCPT2pIadp0YgAequutd
DmY8YOS5J5Ay/g9ywLsVgc0eONg6mCeN1Ju0i1XBZz/Us59QFEbh70FLO+Ron8wA
HbXvDt+lwlwsALM60sJfThMAVZ7eSJ90hc0vU/CxjfHamtoZ0AUC1i6HtvzgVs6t
L16KMOQ6mmkYiUPYts6u1PzW/+w8p1lRCNr5YEYkQz2TA+RZgtQgHAx7tdI3dsif
xXJIiF05gYeC9VqbNGmORw0H8hpkyWhJUnF+MzwBmO8KB8ZrvqTGW0YcaRn1vYNQ
gp1Y/ikSaBTrSJFYtVRFrb5f9m7a1wsrbLZguO/ZsGvXRcWFjXoT9JfCX9fTYvV0
a5QgmvErN8ryL/ePhJqaPGm/BWR0Z+CWq4ZF5Lu8JY8zYT5oBEn+mDAsW4odLoAv
rIi7A59OgaJsVgk7L4h6LrE9pyqykZ+pvxNpjah9pkwpd75FdCIGOQqAHuZlq648
hS+cseFz9Ep96UlNoOzOFzyjVOoOTaM3R0HqUc1d6uFOnFqrwXL28KrxcbsXaLSY
4NJxyrRA2b7mIBE5exg3KWSkNAG0m5XucgbIgceZV9AI2vDOsbHaawVlAk4gYyLc
mpTK7K8upq8s/TN8jhpxxwZ24Z0LbrjBZL3ii70ouvZ7aWebdueB/TPNUAnZzboO
4toJ3FEvA85oKDVQ4KaEE8SkVrZEa0t49sD/ING9e6hYs+HNDNiN56o/jhoZ0zFU
yU8PKw8Uymju/36VBpDitU1Bko57Thi0BOoWGk+pyZXdcaPCOT625aI9BuoMEkHI
l505/97TtMT4JuAAaZILrHgxbG+6a9G7AvFtrIsBzhHQx/cl2xlh3auPgrS3JKSW
g1W8a0cTiTkoG4op19KYRHCCOFjm8skw6zjDD9GdcDV0Os3Ztq2VMe26QckJO+xX
MBmzwT8lNDN7OY8St/vpAxLxcYAnIl22A2Otgvj62xmaw5FW0CJf7D5ZioP2ljZg
oL9q8kTZEH8BKDZ6lOkGuu8bBCOnrwRu7AoT+FSMvkzd20C/nZWRHBvnNtLFSIx5
WFtPW5kx+49KOzNSqY77FWTGsK948tR1WLl64euACXzcvOV7NoDp6RCvPVCRkuur
4iKEY8GOia54vH6SzRBF1s3+tpft5ulG0XpTv/kDcq9UTKM8d4jGMUwf5FagHCTn
0Txw/9P1xAvwOC3Gb5oTOL4fMStPQL6xBw5sKGlY0Q4K9A4hYRy9LqqiSCwOBy53
bC1c2KY69DUV6nsBxOMdqGB7j8lFZVxSMAHP3gOjanndyRCvZwtePqCZAXoSXFGa
pnTYZLLIOBFrH3PXIs+FHI7Ix84YlEEGPJBQ7l5SJjfk7zZE4+twRen8YQi3up45
osLNXi9zzqvpEAzGOV5yOYy0bdVnIj6tIDpD5nZbY5u3qEuAOrL0ZGDyDoJPRFTV
aySqroHvkxld/xC6vzJm3bvvrZ5XplFpSNEH7VGYzYzywDCK1JfDU7ufYYNjCiAo
2jspnXq6Vbd8PtKhzx3seGnebkPz6mlI/ttE4JluPn9SxTS8lShu4M/YH3ANzwji
iMVWyk2UhkT09LtEbx4KLAbd/IFIn59ehzig5j6BIYUF1g62bHT+wOrmTGr6WIxl
8oQsjSGcJV5g81fM2CPgXFq9HoAqiO89rKx8Kp8zFO81SCkGLIgyACGeG4WbhE7Z
5vZIDf+MJCzVxWoAw3dJdDPZuMyo2AH/rTC+cYrlN+DzsQY/9MQRP2VafpKLzulP
PrkUIV/byfkDT9AvevY1dgLzGIECE5OGjJfXqaAg3kNZKRQA00jtBwVZDkksOVgU
U3evh/UoLcY2GMJW0nivGctFzNCOz205EJmpVT7gllgSZiOHVAExKxBwIIlCMCkK
QGHOlb7YpF6xzSh0TVe6draqViHQr3L658WpgLIOcc+w7zfo913sAofsWXgDyA5S
/xNEPrm+mAqJIfb9q2hByo+QbrC9x6UDXGYL/O5ud4tXScY8qnvLND53bmA6Rj2g
VxRTCp0iaooi+qCoSxj+YMx4X8n74aYGrkM5/SqTBEkaVLvq8+N0dIBdPKb5+wrz
F7ptkxQ6rWiTzJnJUvdU/AibfGRZZkPvqxMbdNSsOXq6yittnONXmWjQ1PisytoA
NS8H7obiFVrc/7JFYtG+YjSTjcRN3maDEZ+e2DD6g22tOmSFhGouExKip6TRLtJh
q43LDK5zHhO9daQFbKlyeHxv8lCQIvZD3f/tyU4xcmKfIrvhyZxd/dBDm6keaD13
kNtiZJqzeLxCHKB8KV2zlKaCsPwq1/ZTWNOLQre2HCeElbbgdYP9IoWllATJTZGo
Hp7yMQkZETP3kZzbbmIgUybPFr4KvTxIyNDGqkIoGb31nbsMZoFBXwRoONKvpdhJ
Q9bnL0wO/iRTDepLl/17ySjzWot+ZRamo1LSmmuzGTMSa7B0R9TXU8wjK9AoKtKM
Q9EcaFUgAULSGN8iFbDeNcatZUrCuqU8CNFVJ4T32VlsWk071nl6l0lSGnjwQfCC
zYf+EJmjOz40DtaYEd98DPFXmkP5k2tYPoOtr2SR6D9+EpdJzYobEnBOlPA7aRLJ
Hv0tH+SPahcLTC+T+AOGI/ZIyKdQJrolDbqqYzwIcMjweRRT4Zp1ClDsm1J8pUby
yJUbl18mP+MxxYBgyZiyIGiLimYf5tFEIm4NZzSese/niiv9FcMRGLxPmV4WZQXb
6DvGVKMe6WjLskiGjgNP2HOC1oRrxnFioQlWTyhScxwzPU7TxuPQjmwY9TNYNdyV
pcB5VSVY959ijYtmHAf8kGVMMadzltJABYTrQKrHYUnP8Lo6pg8pi31lyYpYj6RI
5mUS3pu7LoleYrrjWtb5NSkDw1Q34JcoFAZbdx1VbNoVzHd0KcwbWZH/cMw/eKTH
trukpOpFaqZ0w9TJQLlgfnBQNwEBc/NiF78aTAyFX4rukJqnnHNYRMPoLnZTP5Jk
LjCsYvqk8+YDktRXkkHV8xpQHMMhfVjqs6SAfYdLo5KZUEmHj/nyxKB8MzDBgKpQ
JVajBnGTGgGtdLJgkuSCvw7a/bYlitiRyglH+cA8UrJI5r41KCc61R0twZjiBtcT
5WlNchWdWn1CMIr9wosHmZaCUjpcUY2FcYdtbADbdBZc5yF09C2CzI9BLNyi8RSq
4/wHB+zdjp70XMivFiOThLjH/ewyjzypiIxtmaNmcZaf0TD7W2+qyT93kXXHiWu8
a65vj5sE+9auJ8dbTsV/Kn9dfRQwHZDD+wgaV/xbxRErg1zDwk3ucTgcKPTW1yee
/doJv+3F7YUdmHZkrhJd7qop26KzzDp2nyYiuesj27WqB8TO7RUJ0MD+4ELML3hx
yWppGzbjRbFN+R/bYAmNRmrFZazrI30n6aJPrf99MjhZmHi9w/ZKyuFVQu/2adS6
QeSme6GdfURaJxAtEUgSXfPtArb3ImjOmQFspWkoR10x9KdIcR4hpAfylEte2I7b
1ZG8KfVwIGyhkndbCSTc02Mzx3GNgpewVloynp9uJOy6J9OGJQ13o0wnNFCiXAgx
ZarJekOxPCO5T6x9DcF7B6XDS1tOEWHDBzP6rgIkpaZRgW81rqofBkfEz1ojHgcy
d+j/unB2eY5nMAcA0VPKpVGelYEjjiL3HoqYhyZw9GZdqOzTuqc5sFFLO9rPQeHz
wEvVHVYC9JVt764Hns4KuUVB5nE9q/6+1zMYY4zbPQMyjAJJTbOkM0ZzKhNvwLsA
9XcuOm9jMLpzJpuGWE9VuEOyTodicgAJZTUyNyXHXVvUzRoqAdFAT+CIM8yH+Sxx
YP0jkxWhZEK1J//Kfc7m3PKiUsEt5a3mBuOKu9rhqkAxC6pILXcQ24kLPMoSaCVb
B1pvcLY7rhSOG3ggxmtt4jgGQehGVGtui+lT8GyHhcL5uzjAB15jD/LSUUWdLfBH
PSEstGgDk3yjjRj6m/eBIw2qtxJ6csKlfXrkRXEGV130D6z1J5xCRRRp+v9U/zbT
yMxVI79enV12O1Peh6CJdgE46k+TC4iHe3LcnN1DcTD5UpGalvHGxZT0KWrouZHK
+W3EDsjr/n1Bddennu87ed49KqCyUoHyiCaGv3SNamb3ewgMpwl9XRAzFu/Olt8X
aXKwkJlczvUfYujHdPwcZ8efEmaQ+hcetxTltkpuKPrXka2ExDq4ARfhehKdQTXr
+3ym+0+T3kNEYgDHBwVqkDNVc60qtzTWWGd23VQp4Ce/fbkC6T5vkpQ2LMjgrGHi
DC+xn2kIgZIy9b8fIyW4uJ98QfR9psBMwo8cz/E+2zsjyXLfY6vgapksZbdUrdco
/O0rQmmGypKRtRUrhXmJxsjxZAJspavk0NQ4xTNthnjqpgu9bA57fN+n+Ar4axVU
ngUVD64BA8+dByM0/dHtfGK2nn3e+aggQgWnE+83F8jA6RYhsYWLhAPLhn1y/+vX
echNNZG8pzzhq3Mgzx4+B2BkA5CB/Wexh38w8Mf7u5KY+Pnx/7cIxZbyNlHhn6Ls
mJRSX4zxZ4ZR9ZnRzkfSQnx9GnzMAARun8R8NqtvDiJTVhznkWU02odHl/O2mgdH
vEVi5xekZ8JvcW54/FQazD28xXT9pjCMK4gjoUxljF4URBTFhK6PYFyDSwUwArtn
V9Ao9AsEKSUNEywrjO5RiRUG1uXO37zfWdmL5SrLDwU3VmWD4qeqe7IsLbdb4AeH
WgPj+xKosltwDL6lsYeavXzX1xJ3/n0coVFLX2iXHCIsSKXwxPRhn86ICMFjlF6J
mATm2HkUQ/Ms3z8l3MzoAVqXVNCPgXCImuAyreN8wOx7xVUYbJ7fa3YJhq+J9Hms
ddY2+rS+v9DQ0Zuirf5pu/amb9yzDTB0+c7fw4ABOkOMNa9SpFptoqz3EV/WoPb/
O4rU3oiRtlGt07Di+DuRJEo8D9VwF4Np49v5SOcnQeiKOwPNh2evglWdgyYWqYlH
0p5WuhgZldp1EkhUeTwgIPc3ZTTxQT4lo/jkObk0tSnIxda+E1gE2VGgZDWgBaH0
xop0h78DhiqtwjvneQGv3R+Vh1xj75jKEKwxaUAYAUaV5AWtWEedMShR/MZC4JMj
dEr56Gp4CZCJSUMYt4Jjh7M0mZhbar7rk9nME/aEYN0dGPIQLi1rZ0Bsn44aFXkx
ulftQZiaODBENkVjx/nQMjHuuiEUcwG6BlD0GsyGdYIZ5JDJBuLkMEWRifwaDGOY
KLi+Ob13WPXirEX1Zp7NVNWPrGf3lYuwLZoL8HRFkpl8PYIMucHWVfdpipLuD21K
R2ZXWUUObd+w1c+q2UlgB/4veeWGOs4ueu4e7e/4ah0rrlJGI/AJFdvSuXET65Fb
Tr34Kym5dGshBwSJdHb30g3dhlkNDMif0LrBJXyIsyH1++okXMwQJbbkkLxZJKAI
te5Ld9SZ2nBBjzzYCJfWG0TX9jViAdcjMlpUmkpmTRrMuIifZ2jU/31P3ih3GCEK
WLnjETNiD3ErJB94KwxPLefLFZPAwiRoKAZLMXcWPkMUOepMjd2AH4yCicblf+zH
MXFzQnnwlYVm7tq7e6Apl6VP1ouQIiWDh4LScokcBzHfkF4jlwQm85UjXyjX1qZm
GQ+8UTFW4BCU50efeazZ+1o3Ibbge+p2IyXMHKJUbu3Vt588pOcURyazmkb20OGB
Qz/1+gYasGip02TYB0t5Zw2AHLvg2WKXpR1ggB7rjGhlsbWXlI5HhJTzs9lj5Bvc
d2XQDdKY2OWC557Ky2gSZyCQYC6rDrtVn76WL2FUg2wJdtjutNV5/DqgyU/3JIDl
3trI+ZOqf4VXjD1xnRIQI6LVfrypFdQSmGnNzGBer4Cd7XKsMxLfJ0uzyzLhvi4W
VuY3F72QRvGrq2edLVcxPFqZ7eSbbv14Nu4RRGS3trtoMMcRiFYqbxMDstAES0k/
9H937YK/D4eR3/Ie38l0Jcl3gSYC8YtS43ckRa9ud+R9ycuuQ0vZpCEl6jTUiUYX
PUfqCY/EpKkc4jcffXrQQNMY8fptbHF8O4bLA8gDHV6IZSIz1DnEOUvSfvebKvOs
CcGEDRnbS8U6t9bJUfqEz0tGPIMdKy4exsvQSwwOvHn9pSlMInmzgnMXwLEwEfbF
QKf+OWeZyuZvfiNI22yNdPqqJNzAdhXtHRGt+uVx7FUapD+CAe/2btVD/PtPJMUP
J+OgLxVEtbF6KNmvnzKWa6I4eA08tOCwXC10VgQmBI2Z66fv76v7RYSWKQAyc/AL
XimzvTFxNRiSZqgP3hw4wiCngAUpFQ6uicJA3b0bGapek+CNR8o/dYD0QLdtz71K
S3sYQ7NFvsr7K7wXSv7Y3bkF1mj+cp70wnPde+J6rMJI4wQVDo+sJP4+sYFmTCIF
M1DGv2DGlUTNr3eEi10YA6OHijYxlcGO6RFkgsNiIsjAdbVBkioZCBnaOcIdJC0C
V5LwzSNNOT0tMM6SGT6TPW1hFaWL2ShtFZtIYlal7MSpCbZqmLMvaR3p3QLETZyX
19m4qa9dgTBeJw1m1Fy/AC0I2zulZ61OafQNaTjSOeIMIiigo4j5mRrA+2VaC3xB
+cZm80EFRHnq/EbqfKz2lH6YJtvROeFEXd7Rb9QUgQvbbzYf7k9XsbtU7EQpTPf3
vg2RzFn/QhfAZrxdbTF628N5koWxLhZqB9MOLMIIJ5qA5cUCbeim+F04SNV7g7Um
j+i/SKFimekMOOOl6sN6h4tN+yTlaojvBgbdQ+ymybjYHB60W4P0mWfW7gNqHrlp
BL7DGxKI7TAuYv6hu+OEaoioKXL1//fFUghEXcEY0TOCTDnIDEsBaR7K6jLOQ9s9
JcR7r7t09qgIPIkE70pUSuoYT7Es4HFXgSkAngbtoAntj/oSWh6f/dGGWuyJ7wZR
WtscBJgg0pHHwc2kLlAx1qA86ANNQIj9UbpCP60Hym/DMF0XNud47eI97KWLtoDV
wXE3Kj/JhofJuEguby4lwViaEyCbuqSQ7AjiUriZk0As0OI7Dq61LFb2bXsp0V1n
yJgGTf7isgpeKE7JntOPPIBcMRaqk9vCibZYrhHDs9k0KjXP0Ime8j3fLwlyxErf
1SpRiSxh3SDNIJcIzoCYlDwiHfcnXjEj8gimL/ajZmgC0A7iIsKOkOv+czaaHNK+
y0wdvBx72iqhKyPFnzZyhQl8RXLmXw19IjVuGRe9kDmWRVo0DBXCvVdlssPKhYzH
NyByGOO0YZfNGBBf+u0XIdYF1c6ytQ+qdOuTDlD7RKE9ZzKaHh6fGtcsoE0De4f0
VYcHAUUWInthtpwIY+2eI5QAYaszOsGx2gx5rHCpmlx9dDHPXC2yvmpdaH+T1K+t
P9sn6buVosiWrzcFsvHt6n73BHbswBQe8Ji7OYZBXBX4DRzh+Rqc92FTR4JOqWTp
Z4dl/VaF+3rl6WIMZluy2X6uMP20KaW3gFioDwCOIlXLhaokGxpvJuJ9aupBPqdP
D5p09Q90HXgADmrYc7k8fyUsWmfvIqjdqdy+YWEiPSCNddwn0pDpTeaocUultXdK
iNc/Xy/gy+yPUvbduTKD50kSGMonCklNeWUzpbZZZhp8Jh9/q9vVq4iWxbyfD6Ij
fLQBPnyG8FZb6sW/IZeZgcPUHCMj36kSfSL89FVQOtJY+F7SXX2UfPM7lwd+s1KI
ql1h0YuZGVTo47ulFChDNsHag+bYcrEqCwQJT/ri7sYGtrX9oWwstr4zOiMvdps9
HvgtSVQVoikK6PQnKcn/8JKehnsXJ88vl9kIl0OKYfNFqPrx567XcnzlWntjwDcb
8VbmHs3tLil6teajCeZe/U54Ugw8IDSiyu+fUOWhtn259spxG8ujEYQtYEQlVp0n
wRWdfZlBfD7aoL+ftECr1PtIgjM/cgVdU0BB49+inXshI3Hqq2MwtjVB3fAVuPT4
d3BCCqbMy4JajCIuvbddlmelCdwoT4icOZ7Bb5QwPFA2MXnq9SiLO64IwgBACND2
dIbqGfXuNLqTJhjLPuBo2sXmn21nzFwcIGt8lIWuGmLrcU72jnCI1hOJJj4QRiE7
d89NvRlYcUPLKb/eupia2vx5oFz5NfiKQLux3oNk6RryzgITTeK1xLr+XyTp/sBs
7CQbXIvVH39H4TbY8a+j4Dic7LotsjGGAyu52iZj9RDkBx54jPrR28wa2bQrI3lT
tno6v8Pa4wnZxH6fF2oHa+Ne2PEmf43s8WRbi/5kvU3gwo6Gn72HrMvD0TPtDruv
GjjqLnzhu7CodBOFE/mCpmyhuHdkjXFCv+jp0unEs/OizQHbdbXRxqDmS+B40sH4
o4tzK+r7pcTECxCJLryogBRbFRLt1o+74JTquzaouu4ghEPJb66zH5TrPQZ4e8ma
Nl0gaMUXU8VvPqVCVlj0BFVKUPsKYVMmRFdU0MGhIHARQwiJbLzae3j7coq5WvfY
oav1VjOEiFLgKbMTeL4BdiKkJV1TmxrDbc5DM2EfBxMeyGecJ9mcM+TfZe6ZPmy5
o1jn7ZZWCIexHI/m2nBQHrLioEbfXxrt+x+wsiRJuIT9pg8BVhk1QVFnD651fV4+
PEagsgUaybPKrDdQvUOkqvqjGKo83FI3nSUoFW+wVgGtJBVp9EBXpErmewV434Q6
hVOwy4jXMf4OPnWwu0uOWU+jxW4vqEBEVeDY9Sgs2HOdIIq661TkSX3xIkgm+MYv
i76zCRg4Oj81QLlcdhP/TUJxlF85JjK1mDj4h2AGM+GTrPT/T64KCQnF3utTYhVo
ZEVI/9qgOwioZGJX7Ak1wmUrQOrL3S3CHGyzL0ZsMx+YL/VVHDS7aTqoNYWDGzaw
UTd7fqtgwgqb0GGs4gu563+ApYsxdogMn88pHVMb1ralUjatwSojTeZZTd7OpU53
SWRyowlWleW5fpgiXLt7J5UdBUFfnSvYs4fYUHB/tSKjX92fofNN3Y7IxwmysBUe
YyYfCW51nepPXRV1V9eMk8fzbutU9aZ7wVJJmocdQTxka8yVmWId59VqovByW6Bh
7Ae7WuISIqxEDM0Il+T+18EGU8gzzdpXoTHhHseDZHcLGF1+BokrVnAiZAO36Rx5
jaJHtMINhP1aQpnp9ilmnmMOMe+TWgPspnohPmjTfsDguYnpmj8qD4T2L7puSggm
`pragma protect end_protected

`endif // `ifndef _VPR_MEM_TYPED_SV_


