//----------------------------------------------------------------------
/**
 * @file vf_mba_env.sv
 * @brief Defines VF MBA environment class.
 */
/*
 * Copyright (C) 2009-2016 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_MBA_ENV_SV_
`define _VF_MBA_ENV_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
kwbmrgRu7J6CcmJI96XiXuFe0UHXJx07eb/QIQNsxJNwffeC9d8Fc51a65mMaT07
QbweIWTrUnurLGw13X61ou6QqR6Wu9PMUivUwXhYCZZX+kTj7CL8WmmUCQKmxA3n
8sElVDL8brQDrLfgRzVq/ohKVX18o+2JYqEx1eghZeBExbVsWDkVer9JLt89qLI0
tYY4GBOeexJtLu/mYJNaz4Ed4m5DlrEbSP8J6Gp3WC/VXUvk9HPCaVp9Pn07KX4E
6XfJhELaQ63I+OxwHHJnls2zK1+52zeT1zlWotj9QhO2P4wL0s0DECkCIsb29p5m
olu/M2hyjOJyh7BDCtYfgw==
`pragma protect data_block
4iffBB5o+X5ehRtrT5K5n88Qn6QvHvG2okYmAcabA1t6KjNrT5tSFzXCNBWn/AJN
k/o/WPwUusGTpXqPAr4ii4K0yI12bpmwlhVNv1LBS9iUBY6t1Unkt9o7NdLEOXNP
5qy5Dqm6CFHvSTX3s7Hb6N21N6CHGDsrAULHnQxLHLir2O0cCMKJxWJBWTeSQncf
7VhV36NddD8zBwQHSv+vB/nKNbS6k6q8j01zslAPmbcGDksxzNpkQbZWGZIkpqap
7YHOWWFt2aRuGb1NnaoTP0Zei9497B3Ls+KUEog56VmuKeDO/mleQJQwbq5HWiDl
jPfil6xDL2mhMT+9ypmy3CcB+65r/z02R/ErsxKKUE9mmqfNgRHTjgw0EpIW7Mvr
vQz9BlaFWEQFFazAJKObgX1oODmom1G1ffYuOUUQ5UD1yOnGPkgmhicu14trINcu
5GUJnyeSqV2t9q93ncb/1pEgr/Tc839nFhbEBpLD1fOEGaLjc7VmrKPZrqm6DxpH
/coK9NtygqYteZvPktrC46e7pOq80zPCHjos+OBrc2Y4w8TTfc+8nELHMqjxqrYI
xL7TD1dcxIYEkKPRN4unGUqtI8zXFfwawuM7OfPK+LEtSub/SAy2Jq6WW26bxmt6
cynscISXyWohm1VwbkZ2ImAmxgP2dXo2bVvL5F6evDIb/01wBFSp/yQDxpFuzrIZ
ZyDBY1ngwpntwUGk17dNlAGLt6jyp2RfWtorSg6I89P6syxSzGg+IcWTpA4sFDVN
CJINa6nWrMteTw0azfo32mfgcRaVjoHGM/1fj0UnCFHHjBIGcnc/XqE/cEjgI4FS
HFsBxORZoMe36nWVhFRoK/vOlHi5NjYE15I5tiIQWUl+jKoeWo+NUtvfk1gzXfcL
p7Y735aDPqWCk2W2O19AUJb7NK3wJU3lcYLwpHsFv2SRLS1BWUfGGsh8gpN77lGF
1Hcpps2aY3QAJJPTA19FXAUFEiyHZlE85exyNZZp5AscvHZsLPwW/Ersu8/bfeCX
jNc3iQC1PYAKmcfzXm8Sp0vBwjaZG0d/0ZNdL7+fwyNFEp2vkwQFnoT5BWkorfeP
NIz1qDKwl6z6hvHP3xq3b+lFhl5hH1VbWDbeKgZd8dcY6pWsFx7XugDH95ugGSb2
U5iNtOvJVz4VU2OZGr80OqOBPqfIqDEaieLV4+1FYr5xOYec6eftYERpKUCmKmrW
pPaFYIQDTfZJm9sx0VyJmSISNBjuK7w3tZw30iui0VYS/CNHT8DCbflQS30KoIjf
z/nrYtQkC4Jp4aEccX+Uhs08Y6I8ZO1JNCHP1pGlxA1JeSNKTq1z2aX9O0sm7KKK
eUH+K50RXH+sbiT4osBy1WcHUQjsgIoYw1JUOSGqJ4CE2GdGQbM4+Fq6xnZpD0uR
RGgs0C8bhJm38pdg+PSJaspzqqEHPnJeM5gB83H1OS2WzxNCs0O0Ru60IVpvrG5m
uPwDv1kIW9NFyBCHDAQ/0fAoM6JG/25hp55GmDZEkzapebqg3zv6672wiwmkVTx5
jtJC46M8RwjryAKSfpFfBt40RGLTnfaqntcavc77AYhBEE77clIqhlMF9X177ucg
tkR9XNwZxnkyvRu4kpsiyAqvTO8qNRsjJok7d9UVuzsKxUezKuDLP7jbYUAjgwNd
Q1WMW7qvfAP+hqVjFyc+AkX82gGYZ9eaAY3FTLAkD4Wm6QaJRlr1te9MPoMldhE5
jECF5ox8ZnKo/usPKiqg4AYFDJBSGmXydYX3r5GiounD7trqMtG6EfxId6IfHEEi
L1OaklkFoiGTA5gNtj+fu9ICg27e/Z0ZvRTNGp1BBSkp4qb/7FU4+AbvtHG4th95
UJ18AZSUxLUZifzbwqcEzZ2elLU/3yMD018TjU8g2kc/IMqXL1SNApHXGHeEMEBx
++XOSnYoCucWQHcM5staS30RaAGrsN4Dq6XAk1S+xwn5njiTFwKBUDR/4pPvYpJT
lYUuyvDXKe+1cAD6C80W8kLQ4ni5BbVsuqi7k7IynNBElmtWePFYl5OsU1gNQMtl
ijEqWiLmjzfXyALHswCg0udeR99jLPQ2EwuBU82AtwQCxqw5H+z7NPaS+YGVvlFV
2O7JUwn1WLLP1P++kLIM9RxSPIwwk6cwVYl/SKOgi5lRciW4mLeGtrbpYNwXUdny
fBmfoV6qJs7+UIb+vBaK4B/QEn4kpY0HI7Uym3nhRS4ZFV6ptCskfeI9x7LXxHWp
txcJ4vCigbWLL4ct9EOCcKWn451O4cT+p8MNdHT77fmUoLMTBzvZBBeyFaCE0pA8
F3seBILuAZa34hmeOz10UJ/61juGk9EOcKvWgxaOMhfsadWqaVbU/TvB+tAxp6mk
wi4iPxFztzE6oS8Jw8WiKNq+hATB2C8hVe1aMXxT6Pp8L1/u9upfWOZRbBcAKv73
I58AakSQR9h9u+rcs9iu8rbKCfNkwe/AnQlkkIk6Qmf2lSt5K7MpVhvRtdH1dIeH
LNIAA6xWZRP1zqqPtlz+n17FAYTmMgZwMnss57k05hX6gon6oKQ6qniWrLGzxbM7
lxDygtL9lSvcv/OZOY3SWXRsDVZ8/xKQihVJDkz8ewWT8gPQzkZoO75c2BOFBBxU
n7zW1bVGwcDpqOYG997ygdqOKb71p++9KHOtdQz4BN09YWAXN34scZUegzza/6H0
++DjdIKhccplS5iz8ctW74OsGLuTISt5LT6y9GwFsg0SKgX/QmdEWTeLWSb8SKc7
mD+2be+Rjm+6H3kIQoRfC6qJ1EhzKuHqQShhil3Bmwt80NZRhTpR5dhlzJ5Expei
ZIHqDMh9R0kw+L70sX4K9UTz+0BVw3CfKEfB/f1RCEHjtkTsT3H9U+uqPOZJ8NxV
AWG1FSnkWeBuCdQmf3F+t+sAt844R45zQFMBMlUrz8+1H0mqqeDeBBZh5UUOASL1
uwhtI+QhmczgYXph88JEfY847F/trgkD3GM8A6a47tFlq08hGTRevqolugqpN7JR
CqEl3AhQDJUECzpEXgTFTkwW8jztBRJrNBRrjCta7IR7lg5lT9F94vB02x6G+YaU
PTjkE9IuLV+r8uvqn64UyKs1szCOJZ9Q06lYFoiRTuMZHLIKBi1GllFB8plTOKmn
GlH0I78Int/sEYsGZNGkE9b3xjHCMsWLYFwh0kKxtuu3hppMlBGWRwNd1GFXN2+8
US+GEuyDyHh1LJkgMa14tncuQevt0eTL0RzpQWpjNmPbTlDiTJ7HNROjmKxh4teB
LkblTEdNGaPFK6TfLU18uB0qj5AnPYV3sb72AwV9/Ny6KUs14N64SQ5EU/Tv2ZwA
cH4P4Mx73X80pzzlQD+qZHQmwbUGB3OGrJI9whiQpcIJeY55QOhZ0S44lQrqZ+VB
aL3inxq82RlWIjMERcas+KiIJzU1BG3s0V/5CXl3hwwQKCyQl14LgYC2guoDxNnt
ZRNt+bKi8xPsyVZOy7xUC0EtniNefEC+FPavV5EHshtNfwQYS5oVvYA+v1hHv7/E
53WADlzoGhu0bk4ufSt4N24O236kqvyke1i4WhyVDtlRFPhbpcXn30h7TVEP9pXJ
JtNkR+ugTsher+d1/Xb+/Y/1U9KG0nRHXUS+P054wA/PDw6fy5c7RRb9rN8yucQ2
sUttrgIyxq07McWbt4xXxtlXVTWoaKYYPuprm6STUP7hU8/HA5nV05ZVtci/JY/L
81BKncdCmO9AaZOrqAdfL0WMI0FYhQnen/PrKRv2o4x04aP1NiYZafKzeRw+RXlv
bOCUYcxMQFqtVIK8By/1jJtXhDj+wgIaTSXvrJ9q+xnOHGPXSpGH/8V782kea3wl
Nftjvr4QI3aKyMyVN5QzIG6OVXVNjCyyDikMFZjrDdIEK6XLY2cROhNZsYEi3/Dz
oOxdV1CN+/0VLgGF17+vhIVycZTFUjF7ooaug+UQMDCHc7ljt29T2UvpkDVNRNXq
tM6XpMJOxjkMp/w0IYA5tHn6wyAUhKHPpRH+FdB0Q1oSs9un+Gs8o+JGh3uIKJkh
vQFdXB6fys7DmWBHJo01eLgeiLkOVh+NXOuNsipnlrAgrEICC8caRAguiPzjXd7f
e//l8m6tvV6sMtOK4sTLiAO/nH17GjAd1AdUw6jVbdMSokyKHQ6Mc9KADmm30Cea
KXF8frQCQl55lw7Ao2vGbdZPJsbwE1TV6gvMQu4CfVObJweoTCi8IFKeRu+Tn5Bo
OSxJfVsXcgEOhzlEMlpPExIDn4tRj1Uf9JISzJ9ABDwvICBAI2X/uX2fQ+FSbIPe
NduyWzhch9J+3hc13W/JpWyszI6nkEkjPdD5IvNQR5goCO8XFXJG+YPGc6STXg9N
S+dV19kFqolmBoP3k0+viHU+sXtyHity2gplmumL3YdcKjtQuseBO+btYINjflrr
4fMJoTBKEndk4ozPAP+oW9s8soRK7vqJBRFmT+LFOPvhjDOCV9erFb2+tbcLD5oH
3AUZHEiU2a/F53mqEs0FrrtvAOKyQtGMUSGb+e0s6AqYmV96f7ocdxY4deN1k72G
C99ej0eBVt/My4V8kFt0v/u2jwld19PLLQZkCseCNaN4v21PeTUXr9Gbym5LQrw9
gAukZ/odmPKE9asQ/AIPKlLjN8oYWbn95JvRO9piNAVd998ALMCRUb3uwqqTT6OS
x0WFMsGeYQUNEN2HrmzYvLhdQuyTGOISC20Upw2AcVcgjRbxjFo6hVbWJJPJBVju
lnRo7IF5ks+HWuyhSogh415IMJYf5jTmbR4n3VyaYPpY80qZFiSXRd54KA9nWz5D
L4dD9GL1l2A1ddmAEx1xtNO+GAcf17hD0uTQq35rMj+RhJd4dRNkqXsIB/qHwgsw
cwprtQGUykjqOO3a9bScX0bv2Fg+r51PyOKE/q0yVotdiaE91TIopS2zsksfDvMO
3cl7+YReIP29byW8vpK+99khqVoOXLApBk6KVTHaWKUZZv3WMp999Lr/BRwOE7JV
5sYBxz0nEsMHUcTwpTMs2Xe3IBaN//VsjzrnrDm0LedAc6/ca8mhtMFhunArknaj
JxEoj7RpAen6+hQUlkVuQ7BGvGuZuuk3XVN6jRgTxV6Lxq7NuFB+kCd1eSu5oP4z
HJEwSYXRUsjFSbDq/zUyLORbBWhKDPG4IWwa4OS4yRHzNwpU1tYWCToM86i0ngRt
RWACntMNV1gYctB7pyniJ5N3bBamB+cOsnCNLJOX8NI8dJK3x7+3H9RNhjjWi6ca
L3SAKuM6QE+otpz+cfHrjkXcT891LVe8bxcWFK5C33p05JGQs+yGOu5f1+CK8SYn
lFkowoMAbtzAoeta9rF1xxIi6wECV3gyodi2Qdbef6Hp9AlMgfxD63N+lyrBz4x3
J8hxAobkTRi22BXWXkSDY5Tp267rau3QCvOw0/RWwC3chYQufGV/h0GK0aUFa2gU
0IhVj1tclVsNDDkMcQFp0EmOD8wA6zOGNmACazHVGYF8HIWZebUQwwCzXYPB6uxV
CXe78oXAEI0iAlWMNsydbFU5uqpHNBCIXN8nNOsyeMWLoVba48gyvfpr1BWDmJ6l
n/YakHIlG3ejvsAOxQ+5MTHmbdelGQt7WGCg3JwTAEt3W8rcvdR9teKTOeu5Eorg
2WZ6GTG8sWyD8yb+jcXEiNyitn2hlQzQIEMcXdgfHH5R9/5Z99NgcCF1gcq3lmH7
/9tU+b6aapEa4IIVD4tgpPqDEspGA878e7CRenmS8spAZDzthiZCqQeig/JlEmZP
rhaS+nC5yxm+83LQ8MhoKJz5BesB6GCfD0KsPOh4QaHCBq0YQxyc3ad9Cp97tn3N
ayGvjduExg+8Xr4rA49frww6OnDldzRJSbA6nR6WbC+TuAl9b0sSesleL227I6eq
y2WMSJtY1YeqHLb/tpmPeTb033NOID2ZWiQk4Qtrkk83OrDiwFlUNkwSMModfp37
GU9mv+A/anddt0x+sPPXK0t76E6ysSJbJOZPi2smSxKlgB+yOaxwHV1iskqvEkZK
wFneGbrHje3KWUJFcKhdQPQct48x51kQtyX+rBtSphDZpm6y7F3sMUTH7jAws+3q
aMxVlP8j7VVvgHiCp5l9moR3RF+VfVOXkjgjlbMZwd2fRhJ4WXMVSHA0Nh12X1+P
tDkM2SN4U+DCBlkLhZ+qY1V0pbUkki8DsMqVrLjjFwbaOhfJEKDk2uIFFKaqJvxn
2unZqKlFYT3CzTmvAzYiSyBV2JOXWXbkzJm8EfGqpXko5wlXtV0Zs7VngD4ACtLw
9UURcbxBMFFsEarcwoSftsjXPRPnISUli4eP1lwYPU212vU04e7R4HkgSiyN/MWs
oMABZLwzm4epvyO6nfcEa+HxsBVKwNqv4zHOEpS2qT2ZKAeicSJtGU/Pe1OlhsUX
fbq6fLy0/bWv9XS9CVOUZbyqGzoPdMgFG+BQhHI9KKNIkQ/fqNizOSCI8k75ovLi
vutAr0NSJ+AYCJMo1L6OPyyOU8I8jSFLzBRsZG2s09l+HJAnZrcFv1E2EGRt9vSa
yqfroz7TW1Ac/MNXZJahUdA7lniCbL7LBOV9JiVBhO8jY2ZkQZTWG51xjdaE4fl+
s6mvBjZIUMQahCBCqcsdj373+7SmXU0GR88J2fq9oVaTedFuah4BFaijm5cb0NJv
A1OYVqc4TGgL36IOq0sJ9LVT6JE70hO4LfK1kyjSDbNdW3J1lSZQQ67A7gRgI0pc
y1/JYNNkb0thphXIXRsyZsloSbZ4W4Np1/vtqbjQOUdNKuUwaFCnSqIytC6r60k9
uNEMBl5mhkqzsiS2K9VVhuRB+Y66Xu8rVbhykQj8C5v3mw/DVIpPHq7UFUe98/8o
kQ5IVRYRyWO0yVJFsZ0moXDjI0365n9LiAmqsdzVE/e1PdZM22ZJP38dVV487WgI
zr6kzDrnX6k8tXKIuSQZ6R6/HdwzFq2GbJAamSQt212TZEOWpQjZmldAcruMQCjv
B4i/nk7hmdU9exkuNYn8KonEyO6K9uuC/vYeAOIQC3U0C4sv7ir7Uar/aEvXcJ2g
oF5HDt/JV9uv0aNpxbbmuBqdvIXIH+EjZws0vhs3W2E=
`pragma protect end_protected

`endif // `ifndef _VF_MBA_ENV_SV_


