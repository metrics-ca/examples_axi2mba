//----------------------------------------------------------------------
/**
 * @file vf_axi_mon.sv
 * @brief Defines VF AXI monitor class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_MON_SV_
`define _VF_AXI_MON_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
arQpOc9hsToWJbP4jY5moDCNoQN8Wmg+F+PrwW6oDApDRIUiCvYDD3tExJphFspE
svcjmcStkH+1ygrLtnKr2yckvxl4Z+vQtXscdCKiIleYUPBDUuKT94uyj4VIfwzh
NvLbzf1VfjDlPClPVh1yI/fYDxPajth4AUWTqm56Z1ODB3i8NvH3GtwIImVOZgl1
f1gv8oca/QeeUsJK1RncAj8OJHBIayFLYcd4dRwmpTBWr0ss3Ow6sYRISu7T17Z3
3nKL5FpGueQveB1GCTjTn+0PjrYo82LR0/BC/AFLcpsY9VW9hAQVbelA9Dzwi8dS
PLHctdDoib2+HSI2r8oPKA==
`pragma protect data_block
0D3tDGL5S+ZJV2yq85P7XXlrnKH04JN4HZF3Q1kW74rIiiWRGWLJQMD6vRio8ifA
rQUdl+krXnZEzc/2VeZKB5VphkBhfrP+P0hFxUhrLqTASt4Qbo/+66phQtAl9Qnc
YZ0FEpLWQclvmkgsOjdiwqKwItwfgLVagw4k2kygNkMo+elYA9bIJNM9IGIxKA0E
BdxNkd2PdiLrXuNmZhqM8HHqIqgN4Th+TE/51/1NN/I8ymnsrD6KaFlXi/msVW0x
41FEBb5eh2OKfUGdoV3KK1zaLQm02UGtSbXaG2pNUyPiVQo0a2BPis5GMD9Jk/da
EFQL9fhtxzU2xYqEn4L1xJlS5TxIyoC379xKmyR4G/AjAFkdoPlkZSghF+m7gdiL
C+Dx3vgE1QK1XV9uRKrQ89spQG4e8DaNAeso4m2tvG9/TruOnNrYdvKtvpG05uJQ
v8lMkt+Z/AI4E5xveaZJCqLZy/7owBq5tZUzcJKhe9I5jUgJRPcwPDlRFx2KQDRu
wmccNIv/T933Bq0t9UVAEEs4VMEzHl6y4AzqX8rs7BVh67z+k98424AFgvafjh8r
PbifdF7oTVu1fuB83q0ZAXn8oYBuHZ4wL/5pv5rOeN1T6FkgBbFs6O0sQafvb73a
h93ky7Y7olSUm+esccpWMaqkXMxnEo+yrqKVsnxlC9gwgT+RcSjxGUmGCipD+RPO
Ri2bvoFWbZKg3RYd70ua19E5iBmwHX1ok/s9N05aabL6d8Hw5iBZctxExWcE+7TK
FzKn2J3WQieeXpYfST+PkE/98EUgF222Htmf+V4+FcBLyfsVBGw7dzyxL4mWPLHf
MlRlEmRLzUKEiGFEviG1u5BEJ0CGP7G2mwSTe632emZOCSIIxtmJD0Dw6Z8oYP+I
s+it0+729c3JxVEgG8fyc0TLyjmPHOEdIMUMTYKvo+VEMXxenPwYhPaTNmpVmJbp
290jNt2jGgxt5NToFPsQfj+g0+LITSDkyJgFE9ce5KeyrYYOc7VYp/23w48q2MfA
kBjscTcaf+Fyv0PQ2kQlzv0ZtHwWtRy2h0umwSsqo/3tYPjChyVWDVPAB1M7tRNT
BTHKEcrTWj95Nxgum17KJtzBqdpoWlzagFFzFVcrvzr+1BGSmjC0SR6aGZwAHEbL
PRPOhZbUVQgtjp3QwkxA+g8xHPjqjuy5TAYZ1eXuUoUwC7alun/xLZh9QUEbrPZM
sAW9RPOLE1hZuwl/nARsz9e5bSPpkcMDoGkMnwF+3hqJkaUWRkh1nZAq+FYpgfU4
TJ+xaQW/L1AAQrFDcQAu3MXNRD8KO1//jCzkpPMbozO/39i5+UUGlNWBRO3ZxLCv
wL9+4/pjKXqJdHrXffqAoXUO0BUWFXd1rzTN4lVz5Sujzy5kb6t7SfMaR/en/60i
xk6HfveJ0p8fi1rdAN3/fd53A2f5PwLxyMcaJLlqv5oNlx9EogBHdutF6DqSOpbZ
KkrbQoIoFXBFzFcdt6OLajcZzStQfxL99PwMs9VUpdTn0AFyPylvb+RIVrROXgEi
BQmGu+gzVXli12YiKv4S6dccp0ejiRkdvQ8OwmF+PqZc/fhze1QvOtOfh+Z+865/
Dqa1mIsdK0vZ7dBEZHyq5zhRnpPu0ZMMGCiQ+/xTFqw5Tu7famJbHdVi2BNIvRbp
gUIWiEDuVxsSQv/Acsx9gUJ+QXG795qtx9pThqDslTIqOu4D5+gLFYxaOONVcoGQ
jsQlCTXQGfBjuulDbHJibIz3Te95zTA3aH4FirSKhIhJMrFlYhOPjvqAeL2c+LDG
cYNNtyPG+enJSU0bmknWt++TIY7FkTrUK2OjWVhob0VrCIQ/so1s46nnvJS0OalL
/ze5aH8Alnvxcq6yTQAjAk5bVuyZGnZJLqlpLmY88OjkKYywsRPlpL+rlq82UtFf
0vdFRQvO4jpNGkjsjZw14XbkyNzdSXlqv+QMQdH77j6a9SGWCQCD3kRORaDWIoMU
wdf81qBa0dAqWz4l50gN9Fh5igJu/TJ3IBhf1XT2yqX3fjK99+aV7pQDOyJi28OV
+UgwvkUhGphSc42+K+GURA9bujhlYqYcoUBLj0BGn25QpVbG0DmYuS+vh2FuTbKD
NsFsyyUHgV1SYo71SEv7CrxwpXLslfI/9iD3dk8awWfJVekJ7UscDIhGYABDxJEa
Dn1PgaiOM4ZxguUXeIkRuRy9A9by7n09UmmJxplfcteGDdRI9Pu6GmHz369l+tdq
NiblDgax9KVhZMsNQChqow0ajPNDAFJDvg+ZSzoo97DMmQW2bOeJFEQtnZyDewFr
8qljghlKSxG0kEIpkaHyTp7vbdfUcn2T9mHELdSkvWbkDuuZQx+PNd0sizqg/tvG
86EogmX2O2hkmUlEFEjJo/j4GwoLrso/Nj6k87JJhmj/rBT912wTqvIdK4z/DWLW
Ci5IqW1y7tgrRwnvYcXXsUUOCD7VqRPh9lZMYPtL3V9f6j1SGnff5zeEs7aZUrB8
5OxZRxkXgiZIZus5IJF5li0CAMbM4Y8O3KujmsWvSkmEax4TIE/TJ9iWBkEoax3H
UbC36XymDaYg/+mBpTmNCqa7DGfQriM/DYK2E0o+QSjX4+E5JeBhWyVUuCTzbX4T
oJZ33D0UouXHg1iTZuPWEac/9WEn/j4GwHiezFcJM6cUdml5ZO2B4OeDcfd9uyRn
ewA6K/lVO5gUgjionKNsnohpdowSR5aA0DTzTg/PBtsZRiIKbOerixOlVR2lmycv
zQsE2zqR8dfv1twXGPI6yK058ewLQZsDRU7MXQEdyyuNbkQRLDX+hxjSIIJuYyKY
eCgLdEQrouH5XpVc1MfuzfZkAdztU050AzY4i3HPlp4x0zCmWLV6L06GiwF/N7iD
QXe/hzXl7LQpaD1M+CuEBjzwjxOizfWNOMikvSJOX99Pbb7ijzYcvYXcuI4SO4v4
0CJWPUtXYnzmOPPWdRJbVNPhpb9eGRRwbha7ZUHTNEw8IS1dp3usUzAhhja1b0pa
MWsO72QqCiTMyEY7NWSyIkLo+AbG4QGY2WxmT4dqQynCFkfw1isbnP5bbFPbRYbI
Yu3fAMqUBLCucfymVogdVN2uEvChmF5uotCcNM7Zwox9ycwfLsHiJXartc0+B+Mo
4QgIgmiOfeRAp7cayl7DyrtmAdk9nRVtIvok5K8ycYdgzlSpDR7z1NqybE88hdxv
6vBA8XnjbKqd/vFIcAwFJdWb2D5O1BUa5y6RxTfaS/ci+5n4ZcYteiHnn6p6snja
lbhiG0riSU2Udvp2bhALuBqlkwMjzKaia2YB/TNOLWd1wKy+LP5Ba6wZN3fEmkkm
1aja3GdVwLxJ04SlAsuTINV+wK8ldvlRW7J6NgNKmPtj/a9t5Oc15yjggNddjXSs
p0Z/ig1yIoIzvxXrKOWrZQZyswpnalBXxx9X2nvJ0dZL8wrBrRtXr5rLme2TwFVl
dzMJfhl3MQ6o8KDW7+RNhWfMXmpMDCQidIRb+jeEpJRD25AqFuGdiIK+t3s0cn27
LTOBodPWCqIJ2hity0e8WNo9dS9/he+hfOgl1vOAENt8w0Vpa2A0VcUs7My/T2rd
7XZwylq2po32EKWhiT+4Hbj5Hw24EMSOALsZntqbBNRPr59bGk/9wm7dKT5hEu8h
ZB3/ARKGGQDqBtRtliCTRvWA9Jwb7a3AcoMBQT+uWV/0KzlVNKRWlkzSqv5et+As
ngkj69jdAkPjyPerOy3QyqX648pvckctjTw58P0OrsGX5wsQvMBbVWbSFY0Wml3n
oq1LblTxOZFNrdBFWCDBviiEnIS+ksCwXS2cMHBQbBXW0lrCNBwmxMzJclCXJmi9
hoGbJpM2zK220lDJbVV90WOrNR0PuUo8Al3+B2/HoB2dMr39AvKZkIKSBslhuhUT
DLR5KKSI+2svJOeonVcjrZdy8kzLHPjTYNQqxGKmR7TNk3eyR5dsDgXMH/en2/l/
5OlTJ/T1FLChAVs1CMl2YQ7r/tEGirc6pnOWHSKSVF8JHndq8vxxY48Zkg1POxDK
LtSlJUgHuJGYCv8EhZwYaoPOVmJonbW93rXNhlDlMDiAnUk+TtRaP0rT9y6egGcZ
ljk56NjGbp7QwBL8F+kFWxB0Mgf4BYKjwg0o7x85VS78nB22Gf8yLPaXCUYtDe+a
KlnohZIyJJcsN5d7o+ieG9tdj/M7ZymPbYOXGnHhCEtu3Z4ssm0Ad4DIGdkOsieA
0rEfxUZJ91yuYrXnbYmLWa8fobR8mTNRp86FYEbKbDOhZd+CzUwtDJggHGHbK6L9
eKfX4QUi91ZkTIVHxRfwFNpS9Vj3GMYNBpAclmQjMFZoVY2GobPMZfqhVXakYTCh
V3A5cGc+VEK79LDBzhITEuF1D2FIw8e49E5w8yCknQUg3JaXvpg6fBDGGowS7sf4
cDozeIA5Z5mpNSM+8fLYQzVzVtvNFprpGB/Fi/aAJfmpZtxTqnXW3THBpbOlouAR
BakZGNqhzyES+LkmUT93OFxtFDGKu6Tac6By62UEFjb478JOGZT1ZbKkF6hyBYuV
ZfU+OdqmDIr0VKAOqqWbAPj5UBqLHIBaan1lHFiOd76cniedHd2TXoXYkNuxqTP2
hXpxIZ9YtyNEKRgTazWah+47xakNPe6Tz+b5yk41Ma1kRNYwe6bdot4nQ1rF+y94
e8HlqQHJhOej8bMaWkoeAXBhX7RANVsdPdF5htXKtR0xedKA4dISnmMqIq9xiaoQ
RcMQUC9Sml5VRt0ELPENlvqHhBrPiwCSdHlfrBh4YR5Ur4XE2sw+E8L8EWPVguDw
n/e7Nmj7/1a+onDkIpDo9z4rzyCQvm4+btltUKzc12izHAIPbiuALtv1yBkEWEW7
3Px/Oi03TO5wrne+emZ0RXalF8zywZ8z6nCqBiHAbiP5ty/T7HkGW6PwnkljE//u
2a+YL0azJiN+LhzLQUvH9Vcq2+ihieBltINYMUpJHvjfo37fgo9+1C0dMFf1qHTS
E+r+RjJMQ4F5zyuAZHigWSXKNTfiMfvo9HA4eVROg4IVHKNEse+zDUpfNPT1M8sQ
nwL8R7Tz2T/+m94jqwSzV1TF4Dql3fH/tvVZdZAxkSVseV4u/iT/otYKxW7BckuX
jArT9z21B9Wj5jg8DayTE/uL+727FgyeWmSmzCLWJb3t7ZRjWYE7nJkmN4QocqjA
0Aur//t+tgm2QPvivP3AuBBXevvoZbM0c67X5O8h2Y+y/vsGPPuvynAngrkrZjbJ
LdxQuNzXjCSKoEp7nyt6dRxK6gOhovZon3LPlgiwkZDrltZ+au+dZbqnAj5X8gjS
GvDIgfoi7L7bWz2q2sMMHDytaDlK2Jj3RFyJrfmEj7Q5LUKrOPgKOkKiiLSgC0+q
SNdmN5NjYA31l6wLu1lBG5AzcVnG0QwicoVOcK/uOj1YMBuQ2GWxoCzK/ncFCe1Y
yEkcO0gJFFqy196zHKXdyPsEap4ZQZkSStWA+o/w+syYlhEHYjdh9bLLCqifNwB6
jRxPqS2c7Su43+jlzCAH7fotLBlueSwFEOLcGZHcRyq0kxJCRrPJy12Bg5YNLSTY
Ha6IY5OfQntCYzkk1+enl6Z1A3q6937Iuwih/2M+1+FVKFBpOV0DVjbyigDLF3/B
ziyXNkxSb8/1sIpND/fMKD7aesi7V9UIhZEXdvs5A5sXdWSsLv6XIXHm78LwoZtb
faHpxr3D/IlPzVNphjwwcCivREhblWRfdsDbGzgU1RP081hAO+WoYpXal45d0PxO
j2r+bO9d/7R2HGcmkZjLSAsv1x44En6qyK5ixDqe3uXKnbFF28Xi5WhCs2fFZi4+
2uw5aGF0rPsl+pPU1QEm2Tz7KyxtFomZ2+2F7TE8qpDB/rCtCcMAXFEDQ8Nk7bnj
pfLSbrBhJalp1MoYD8+XtJH2fhIraDDIkdOHjmZu0LFlaTFIL9rr+ewKH4lBLGnr
1XPcQzXqrdDsw3KC5rDZFkjWl8lzBYsOsSNRKSAdx94VdzTwhqgguZtJ0Rs0UWlB
I9zGG3JWmGTFY6pruKery27vr4QEahF0XhxoHRoDxhmhUhm0/jhPeiOXuuJPSFCm
A610oOTJrWlMknJ8hhTknLIVUP3noDc8574jHuqSIwBZDUZoQDIrkzkc/0WEYiw7
iYqi7OodFmwchbEAWbKE47ATfVQEJ7CXN6XyJBECtZxVAur4SLQGyRZ2uGDMgItQ
ekxg2FFgCM1RafV7VSQVTGiB7VWPMTdTdCdgSBNByB3yl/VVcRhUw5QIsyVAwU1F
0XrbEg3Ahf4uUK/KzM/wQk2czh0RiFA3iG/FR8TxXacENBbixTsX7WK4Inl6wlcn
5qLntXwYzQB4nBYZepmwQ4yx6irgQzG5kTWzQ0C+xvq9kq0Ovo7Je1EqZ5H0tXy0
mmSu41Uj9uFYs2daE32R41vN66NebgKB4ds4shtNyYagK9j5DUB3+MyeESTzI01D
8Sdr6z1OQZ7yXXREKgtqrHoqvwciDaOFAUemLIisTtGQ0rhalUNXeAGxjUR4opkI
9fx5SUNaNuvL20a+I/LMWte8TpvJSzV2O3odWU4+jnXr0rmSV94ZmM30bMXrw2GS
w8BxIP4av5TVMW3PxzTZ7JRJBJi0/v2A10WE/Y9ddyg9UsAF0epk7JJnMlUEmo4r
JKtdbYemJq47OFwbdTyE6gzwBpi1duCCul3MAdb7mW7DLUFcD6RmgspBUQNCsTOd
N6djppGdMh+t0VGUPtxC/lb7p8z55B90OxrQ8QJJ/8nDjlnVGrJVoINLEg41fx1B
2UlsK014goXHxtVwPOid7oL5MEMkKMsCfp4SLAK7DrRRrD2c49p69oIuZA2CPYPH
u0Aw1VUmdbX9PbgVxO6vzMC26mMgb31YrPFwAyyESpPtCUsTJ33r2CAtCXBbESiX
X1sxkixtnfTAUABzTKMLmmPZMgZczxcZqyBE9dVxfd3nfQD0ARCjo5LjD1+SUaY6
EtVPUlm9PjILScUjj27gpv3cXk1QTMGc5MqHiDTwcDdfxDZu2ACrAmESlZR8coMm
sb6qVQTne299L1Q945kLCpN7DEHxlR30ja1s50ekiVEJ01k3nAoOyCvR9RpNLliE
yi1Z6eJxiRNH9lGI4wXs4KvGRMyvrRCkdg4kT1DqA2R3dGsu+iaSwfBr246vmkEv
0+lh6l06ep+tokZEtZTxTC9lfbMN/j762g9Iq/dPwBkZkNQJOMl1GSWsGUNVB7z+
fvJwzxoO3Tvso7ZIoZ4hqP3yvv5RgLF2HXWLZDdBbOEHVjoqvBLQnZdhQz7dnARK
owgoL2jA7KLYTKgMy5meIae50x/XUL4Gv+A5HcGXkGiYRPoMNHFNKJW8i1KB5mci
pKOL/7se4GzCyhcVMqlvRBMalJK+kck/ne4cHT6g0oWUv/Q6mGllUcaOX7ELqzmR
rtCIScBu9akH6Fs5RAzunVgVvczBjSQq3BMxu+SvrxS57gkUD3hlkeIx9XVPvdQr
goHnwVgu9ZF/j8M3CozCGv4Y3CHOulR9btegBYDGxyJVNmF2a8Wj6/bCmc4Y/6qQ
5ODqxx0eeZNE914pvtRhrvjBU8LExBW6zCuP5XXtAykb5Up/t2kbGla7y3WvHaGX
Qkc3u1Tzn7bw+j58y1pf1LRu6r4QgQrWjuGTpnwvGx1QDb0iMyvzQsogD+FeqncV
4bO6Y0pqRuXsY8aF41NFHbRAQuL9eiAxIhut5Xoz2ZB9AdXDyfRP1qKQb/+XEbrq
ZnH/3XEoels8za2mf+0avnS9ndksPKQDrvx2/6fRvmreLH6KKajzZubUCGCyH/pO
HQLYubNH9STOqR5dxFwJGSmjw4j1yy+fbz82ygj8Lvy1coWRMPDj3ygSC5ddaPZ8
FuPY5DGFgG1/boX/ueHtaaYIgeE1DgbHIQlXth64Obi7hRvqLwUieUGSVxmkpxGo
dLBX/5+vo5qPHQvhARLIXfhJqHc5laejO+lVtHs+iTXl47q1vlprXAkxB5hqTVyG
YwYOprSCwG0QK6a12ygfyoqtyZyYN9ees1Cn/2RK07NFdfIl8TEFoFgIUxIgXccd
DEFvpT3ffL5fGF0+9IxORmsRqifNwfoV/kRUSJ31G/LF/8ox3hu+2tT/igBkuW1p
bQR7CjkaqLBC5zqwQJr0bnewxKAil/ClNPy6P4R8EyKuH4wR+JDeO/1WsEaZGmS6
Oroo2QLGd+clZqrdtptUYFx+EfB/G14f15tGz3QjkBO0SXeJESXUF6Kw8C1Fg19+
GlG/jFTuM8HgKXo3ckBp7FMg9UyVRIXplTv3u064wEADdDc/SEDiIaqQS7O70BuX
1s4vuQGRWy7WZxVnFm3lS9bRBqjSFdzkXbpjevw0u7Q/UQMZj5luQx7oTWQMdrE/
B5BoGv2VW+gecZETq8IOKS8p2Bkyu63VQ7VTikS366eFqBr359JzXu5e0GSRZ7cE
HEqv3ebgkMZuO/Ri6/NSvyjuz3KbKuOTkfuZGdH+eoIHlKHGopdsKEmM7rMP0M2P
U9xc0ulTKhLBH7ft0Y9+rgLYWTW2c3+oc6xv93LHBQeVeWOtfWzxoegyncUNrh7U
TNMOrh7O08ZQw3jvSTl9+K6hGeKF0iCUwV+1+BdYlueQNEmsIMLzmJuJZ9BgzVNi
3aPUD569D8xToVYB8w0OCp7+E6DvVC/MpwaxTglSZnXyv2kZiGpFJg5nrBRNM0XV
eVza7LLT5uzwKlyxNP5k+lStEGSX6E5VobC8xvCc0vVsCPQdG9iCuR/by/+h0QKS
QPbl+1oigOP5JA++F0XM+SpFv+3nK5zrXGjlCvR1ur7Lf3NhSOu+YLY75Szqwo5+
q/+brYVINtUlY66Lg3t5hSs19wTDjUtbM5HHHoaCHjUgkpvJ32vdJ/n/CAxm+Rlh
zHwCPEZqbIPECteI6/u352ROHwMEiosDV0SvID2U+0Xs8nKu6r+mmsHaVtB4SVtP
/apje5GI/5XSiRUeRfbi4JiJdMhGpK/TVKMtUWpzKGLnlVzF7hgBawaQSjo2Uw0X
VWpV2BSRlXk5XDgcGWn53wSD5FIZnatPQwuhmElnCOd+W7rUC6Q1wt5tlBdBXe6Y
SuQOIU60yv8Rqfpu/1UdakvrzAkwvKEEt7YmH9esJO0VLylWSDyr0VtgiF8KyrGn
yI8a7Z3QqYFRqhbL7+X2YFGPpwfdrlUe+2v7ZKaXuJaEawxyAd+RMQz/PNjk9X2d
Phoxoo2/iN8oAcidpdAjrqYE50+oJWhBI6iiCRwVs+NePryCNTECXYMMb8waxghq
MPXgeZEQVELy7hOtStim+F+O4QZd0P8xPFrFp83jTaNNjaWMezYnWWB6qGCVL2fI
urI6XTu2VSI19KE5DEmUWTe6hOG1cVrxN6L3kMKEjozJBPCF+2VZrZ1rqLXnB3M6
2VRKKzC+oRB6btTioFj3ywdwzWP7AN+OKM3DZnyem/Js1QP4ULuhrW+bdq5ZjivZ
lFu04RbzFZYvB4+CQufQTJoFOSjhUoiNK76G+y6VY3QyPYY5pXJy/fRTuJHJ6Ox6
3dZbEjZ0F9wjh5eIffESuEAG0cl21vEA1LnyjXFyZ1pcA1w2eCJB5IGcqMxtBUZ6
7dqAIVMCWvSJtALADRBlEl535w9OcUbU0YZLHc0BuBy6EmJnOcbg4vNxBNfzLhzg
vjeOkpGygcUilFU2H/gVBplN7a0+p1E2ONw3r+dpWb503FnkCSFnHPC8igF3xxoj
Ne9EGp650LBCeKkvqgsJDX29stB+Mpq8BnTWH9B2RT3l2g4DZapJfpTcmXx9CiHb
54tSgBZXpn8J8L6oDInVYuvtg75sLD3F5635MJFXDVbN4MwxQJC/wbJmqLqPbt5J
4HBZORx2rolY52u9kRV9r7+JvNK7N5pnrMaEUchBH1kbF6CjiRCffh0H83vpOGNe
z3NG5FdnIgwaBb/eQAPQ3mi51Bc0Lxpx1FbT7HCV4qYybZl7T4ONnXkdzs4HRkXr
pwmzda85GwUHc9p8Eh/1nORHIFdmETVeM/NlMGnX4n4m/wzXcxNwEGgpqVZPZTMK
BbF3WFTFHJenO01am0dazkRbBKy+WrOiLxowEVCAgpceTdylQ4hx8K4pTMvcDkXT
ASEASXt2ejD2eaKfdRz5nrOay4BVGrPCTwwMawq2whC/Ku+MKqaC1U0/6Th5LZ3E
Vk9yaiYabWZrNKKOEn5U6nyXaQXY7xlq57DRirDlUBzr9YS/nD4HaHoysYM2oAhE
fHg46qLPX2XLiqzK88omefozBYzykY0affNw5YaPT8Z6zSxntnLflMhOuGWKWSL1
9Q2UnACmJHNOUNnI44dgUtRU1S5tsz1N/NNx+/Ibyh6D8fckgeZkAmEtKfCO7pxZ
4viL+mB3rntfV2UPxUikSSSoYsqkbtAetfbTb8GcqNH11bJL9Klf2mKncHBgBCAm
La2KkXRCza4qoY190BT/0gB5KfIxnO3XOug5s/JThOClPytjETZ6Gk7eeId7qqs5
3VCIiNzi99U9tqFHeGAx21EdMyU1OUx3G/O3ljZDXXTvF7pqXgSuq8bPS3XOMQlH
Nzx+ytSGXfLFgd/7e92ufzwj7h1iWWTFdj8Al6Tsc+/1TgRahdYv7Y6QCg1yTgRb
62X8QaFl+DZVQmVt5p3TLxxZStlVJAuTxaq/LSXGaIlUNLRj6sDrffW2UqUBDcIk
gG3ke08d7Ty3SvcZOBBaxrZTU26YFkD21DjnyvUblYQ2Y6f4taLVqZNO8H/Wmfrz
eWA3Pjwe+dhkhKynEZQTEAfe+0rcKCGDKBJeKBS/6QZNrY+vJBbhzWxuGgBhTvkG
WEA4OhNVj5nMN+rFwSMpUYlSOZKgAuUu85ETJ+Ed+R0+7PpwkG0s+ANViqL1eoic
6syhPF2MmS0FnkcmCwfNvwVgOvDNqjaAaHaNo/+SBbrXmd9QXpj669wHnaj0LOWy
0mH8eCauAexlSb74F44cxlcmm8Luhqt/ZFEDY9821k2ceqi6R0w7/5zmCq421s5w
F82X1B2NW4XzDoKwBwN1QIf//hX+Gxe1eBTpj+ZR3yqR8qWfE3/epQS8hfTpsdwJ
FbFezf30JY/vWqpj1jWgmvRtTE5v+Y9EjcWTITXBlgDYs4r+Hl9+hMD8APYhj/9L
Ab+ZMk1QHXBTM5hq1N9I3Hlap5Gl4DWppBig39De5f7rakXVateqw8eaLnK//W4F
qU4ik3dpO2dDa+gV82TtM+DFTYQpTX2j8nKvOQbmw7KqGktc6lSFQCQ/qBW3E7fs
J/VyDzUIzZra3puABWjFpWDVLE5vq0xyEws4I38ZzV3nW6M1nuHEdmrIGnP80Oa1
9H8XclEhjoRoZR0XQYo8hSU26YI4qBYlVL3Af4gZ3HM=
`pragma protect end_protected

`endif // `ifndef _VF_AXI_MON_SV_


