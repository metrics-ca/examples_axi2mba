//----------------------------------------------------------------------
/**
 * @file vsl_mm.sv
 * @brief Defines VSL Memory Manager class.
 *
 * This file contains the following VSL memory manager related classes.
 * - VSL memory manager class
 * - VSL memory region class
 * - VSL memory region queue class
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_MM_SV_
`define _VSL_MM_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
lm0jeLm3DtpSlUTI8qDC+UjD5XYUa7dZ19AlV/GSZQTw98vCbTvfJzPG8lNqjoM9
IiLUyhST5+Bl7DgrLs8ci06oVvcPGRw1UrZef50Z5rdJ0DB3wFebx4omd1jY/+1o
CHaTMWClWfO7NVAv7y/o8ePqmddpB+BpT39FBIiKO66ifI/s1jC/2XdxkwfRhygf
BnbWt3jE7/RI5a92SXfrw12kc1DZRGp0sdlQn8dbsojV5uzb7cWR5ZBeDrD/vPHt
6L1qPWKElJcHEsvy07j6lYYPlCdulZi+fH2kYno0SiHGTZc1uhc6R1p6+t7H6JLh
Ne6NhDBUE28aeQgucYB7+Q==
`pragma protect data_block
tXAK8lOELcM2Q5F7vPozph9g/9qeiq5lzZP13B1FbbQNDvkEpRyATKGzcpo6LsU8
X7XXSCcHCGxQx5QesJTZZOwMOvpQFzRlesY8OGkv2QDpuY5G7Y5cnxENDIfPwMcv
/sNbfLdbm200jJvPRxDqhXRN3RAS/BoymBNPST5KranlqECK/3lgZ+UckrcbZr2+
8gRK3ztNFPODr/0+nadseayi3p2S6SyLwUr7XiiX62yAPWrRCR3eeHeiMHmOAvpv
CoVEaKqE0LYynFlFswmFzS072DplOPa0hwrOHhQgtsjOwplsyarPhbbHXL9syeXx
xAykER6sbIzWjez7YjjZL3JaZHyNGk1mkigzyE/y1B12XIJ7PhWDnG6oE3ZlT/MO
Y4DL93gIYLYePbffHFrb4nQKpdHrSIKAEeOs0JdVC55PLFAK25OmEzOivhS6mjAX
Ck89GFaFf2QcMUPPqAWfXmWKxtd8KBd0mvnC9WpvF2ZRI1vj9QDTEq8vWt9UhMfI
s6/9CChR0WFrW+8Srz5UcPFpFYsKJxG8i8aWv3Or7AKkGQtN6m1FLkjXaHJReL5d
EWccjLD7v40KGkCsNbxGQq9WBgdWV3VcJSXHvtWlRhXLbYSssOyVnERheX0g2VYs
H6sw3g2go+vyXDTVW4R4Sxb0YjGhGm90dHbROIMB1orJfWIMiBjo89GfXQl5tK90
YyTdNBvJxMzolqMsJ3E470j4rtk/1iAkBaIMlOEdL8RAPHj9YsKF/X5o3pka+xjF
SoevzPBaD0zNNb7nXPcmvUzVw+AglOQ2cOWIGBwwA24U5xojKRMNMhb5ozmN7CYj
bB69b6upSyjQ4t6MgTGbyFOMjTYQpL5P7N1lsZQHdePdGujMIjh4O2EE9wyStxGz
g3ZzwvsF/ihpsCee9RoPqobeKFYjbDl2ybM5kXJWHfwhxCrBgPta9X2JORWsWghq
jpDj9t4hSbT81L6D7sOAR8DJeNnSxzFkL0S+p9fBv8ghM0nKOXSQ5uVwFcdg8TOJ
9nQ025RU2lvPi5jlpX/2m3jUEYcuLuB+HQOldyCrKuejyiqavW5pPEjBi505jEz7
y4OuOITMiqia33c98hJyCjgJoqTzvZqc9u2zhiVD7vUZn5MjkOvkeMeEIP4t7Rw0
G+YPF7jOk3e1BOFiNhpaPDxk9b1PVcSM1UtkJZ3kmJTZXQZk6rc3sShIyYygAt6/
2Rf6Px5WRErTXlZXH3P8zTwBApM1HzS+rTrcp163bAytPjQxEmAZ6W21mqmUcKFN
lg71LfT2LJEER2krP1YaVqXsHDL99VI9xnJWZiEtVSD+ULuCCvQbT8t7uL30kvmu
iV3X0dw8j8Hc1FdGRDoWCk9Ixx2EtY//qzlZqYt+Dyy5MV4VirrSf39CuoR5RdMW
tVvX3nHDta426EBw9dGzH4eKViiRAmJqUC3JpfTjJYEv5tNn6sOzCzoiJgUpoY80
0zAx3Oaj0+PrTthe8MNn0MS23EFhePqHnuNcQ725DiralukXqGw24BYR24KqMR8d
UPT/OJqblHnuBJGIhnPwBsxV5vlJeYPdLI/XlnGShNxo+/xnOZgheh0nuvz01/fx
pnGz0unTqg09m1d8lJh7S77rmstT9Ng3ZpRz3mdKZEC+suXfGqrjJpzF2N/RTsF9
s4RFnRzvu2JCI/BeJVt/RBbCZXivcHILNk04ao/HMN95i3rK5wtyrabv3hZEfdSW
oOhB+9d3L9oJgiHhotTb4EBxKtFUqZk5/cKhzUDMDRmu1L414ZsMZdS9mA6eZ19y
wIXpPUTJYe1wmcsBWWLBikqmNP1dh8dkS1RLB+JBy91rG2Q2dZPLfhcDPSRAOd+w
MOFBOLFFklLrzgM4vEdSK6Hff+OZHsah+IhydCCZejyJwC/e6JnkH5beYOL+8iTg
lP4XqeplkbC9e34Hh4xOLI8gGQ+LOOAJiZX79llkoJgmFTiv+YPK3aESAXup2Ijj
BZGWph7L8AeP2teT0OBUj1hAMeizS8SpP4QfYa5isgiSVzutoXUmgVvncAyCe8xD
WIFp3bKBxXylS5AVgICpppB0/Iu+ZN5VI5GGZjRmha6B6EQPmNot/Q8WHf0kaDzv
qa7tidupFuQ0iOXTR4miIBFiRjQRfEoTUTt4vi+snzvjJgrYd35hEORVg8tDS+ex
QD8GxNQcfAO8dKtQRyruq4bbQY26L0MgfoMcWclzn5EHHrLKi936Y/ikFB+yqM/r
1GOQP2WIjcQyuhg3eB6rYlrqlkmeG3nB+rHJEYqNfcdi/Dqfpfv5ZztrIGFhtLaM
RKPqTEjwK2Apk0HcDIl6/I+kwenXNjBMa471W95T+qI40Kxt/heQzAaGlAlrQZrH
s+qSPYqrE2EqLdz9p41hDrLoboPvEwlNSlSonQ8k+ezziamcNc2FHbVFjTDZL+09
ZUbBzHx2ltY5C7bHNEq3+yMZAN7tsxwktMb7ko4ke2/mqPhtYSaBs8QRdJBY35lQ
KnX4775C7j+eraHzrrC2n/PmweDS8lMWol5jxkR3mpEIvfGs7JKYau3h3sYBS1+m
0MlWr9ee3GlMQKho/qj0tR0E7J+fO/POA4EkQODj7IjmUNelyzsgLrYidzttocHS
qeoWzX7YBZ75Z3Gk2+Xd35RQ5ONvA/MTTSrKWxN3D9IxOQ1VGYWFzr6nJIcLZ93m
MKxRoRcriurFStE5e3xR2iDOf3Yao5KwzfTHQ7E2m/PIEbwfB08+cU/c2EZFax0y
K7zS/SSxywsyCKE6OTWgjdXYmfIcyRZWyd0lZXQVrvAOkd77XawPvWkMD0HqUM7+
v3G+Zymw159Sv1/hzjKXBPY3hOvngCjOj5EcrW4/Z27uW5rP6uLVwhDYShFXCSk9
3s4+cnCnHRUAa68Z9vz4i7IAvOkDqJ1MMZmAbzSnBVZqgCbCkRsfG3VH+RcOagNR
RWhXQLukB0AdT4YhlDPy5CU2J1BffxdVw4bIgDFPdMtKJPpZm6mDZRy85bpRzAyw
KEhTjHHpuBu112K+yYGP7sRwwbJYiBgrgDUEGGkPaZiHupnE+RqueuljHN+/Ht/Q
RCVKD/8XhNdZM09eb9oO8Wbyk4o2SPO3uYaRg4+N8Y0DUk2iv0YtjtktEDHM2c4h
v+zwl/cJpMh/iiMVojyf7GQOO+a+VnuQkkEOWhGDOHOyFcY3J2wLI9mr7Da6MHm2
W8wR8LRtuSOigmfXM5KnmDMH8tlpzJ0SCMf+ypTSjW9vEdACo3KKt08cxCR9fHa0
crrgBuL+5VMvsYmMpRohv4ZT/xP/J/KOIB3TtesFnolrRWX11+rPdjzVzCWr4QBb
LSgB6FwQpGJ0ArFK5fFy7VCMwaLAgo+GxIWG51pN6nX9bggdrt0Xz9TPiLKlGIxf
XTjr27IkzBwY9GNKzcMGRFmVQ5uGM+Jx52uAO2XsUO4Nz15Ce90fBnn4fdga0vyG
wp+AxhBD+vIYShBTSpH3NRqZTMYjb3wmXb6u1Oo81kptMrwhc6fze1/caVEBJqoL
VP79bEUpljHT56IFzBZUfVbLmaWhwOyLwZd5xVxleDTcpaxe2sfUkoa7R9G4vd7o
0z3ZaT55oRMQ4kCx0bNzyPGrl98U5WQPkf3DQO+aOrICzx2/4W7JnUBgycrillNI
aN7LYg0fk4+bVP8yj6GDSE77ejNU3eFAj//Q7pkFoy3Q4cxJS0wUc/aCcAzdjOy+
iSYeJ5xJeyC+gKkLAsbKItYj8sp2EvuB32NWhBs/AAiJHTJNUPfLL/pSZjxrl9Bf
LLUHR3Ep8NKRyyN+S00NAez0dxA1Zzzbm4cVFxbJ7QVc5gUyMcFs5vaEEA6B/y9Z
BaY1VaczhNKLr00J8GCFwPFJ4q/3W1RAh29PKn/lmi3Mp8SnwS2tNgLxDfXy/SPh
5mw1NQu92rEBcXj7dIdlqwHPoC2RKWW+RdVnnoHEXrpHb0dV86KOEXY0t6Aj3OvC
ZxRzY0J19NeTMbGvTfRhK2B/NHiKOVI8rlXjeJUmBZRxk4KZ57PZM5cbWn591XtM
o0UXwxMvvux4yXeAlZRU5kV2S7mZgtn8kJ3kDuJXgmCIXb63eRgtfcGuefyqlQEv
z0ddgSQ9eAbMH69h85HYS0PeQ5UA6pB02aIWUF+rPHBg6j3NkBYLD7qXGX2yp9PQ
E3kQq/5yEcRmrERsT6i+zZr8I2Pkqvy3j0qTnRROUkFc+gML1v0orKCLl5tlUVxC
8lmPOdIrUZ4RK4XPqi4UgdCI46zWIwzKqt2bLIwcFvSCBT628w2yt8eSSLeEqUd2
PwPvFpwb7szVG1Ddt3lLD61D7pFp9aVaCdj0FoRJ4OdsQGEITPG07j8Ru1RcNWS4
CjZjd/3FoqJ4PjY2M+CGGxX4fSF09Tcg2jKHY/0hgat7CdJM2AZchB9H/iCQicoD
+kXPj9cd10JbxNiodHavQVqvfkhfjmsrVQbPr+9sGum3FUiQa1GE8XZGd3M4TKN9
/L16KOvG8VXIqZ/to6KAaajJLzVrlw/lhoNocTBKABIz6QchkdeeflB3dCIEbgMN
49XSGgzIvmB4V0naQ3EGEjXreLObCxqaOHh4YZzX7rl2+08QH2ek2tN4oLwyg3XT
TjzprIfd5obepn5tH4LYqYWH5Bma7GsDoevkomY2mgiCGHV5NexUXX/DWwyS47/S
AkjH5/DCZL8KhCHKqjH6utTiTIPAQT/UQ2iiMZZOJlXsPtLN1ouRcsppYwhXvqM9
JQ4rd6Zm82CO/xWzyrvOW+PG61ufWJ6zo53G8SsjFWLYRQvEeO1GJewtPYrqxdPG
uPuKkuRA8gm78yI/vDOczwydUuzWREkubxdg2eN0b7TYK3sbZpHC0vPOngzV7ind
Coro2gqBlpOQYZUonKnp+nz7ZrViZZMO+2/VUZ7YbcA0z0V2Djm/PH4Ww+3BJAVH
b10Tw/RNOJYUZhPLID4LKcrjNNzh/oMRzBV5pwip8bqmCHDpOnpq5km7g1nqcq5R
/gb9HRZ57LGXl2ifZ2vRZ+gE68B//IDlG09xCaSs6smhkzFHG9keI5R3nM4FmUSS
xkTEDoBgDHBrFMXN9rzce/xo2vwYGEqZMo4xy16j7XgQH18d/6YQnUx/8a5oPnAE
ZpBg782+KmfL5rpwm2h+ZzDMyMLOlUx3+11P/n70SBz3nRwRa8kVzvgR2IIW9UIl
21Y22pfq5DJfjt+vVJx8YNl6ZpTzlxlfR2xSYDomssux1lrwtlCbEN5M+oWTnh0f
7R4y/2oNVU79bnWTpTpOvFO79cFRh4HcZqmzb2SsSPKQ9/AUVyVMFMkZle2WIffy
fHeR2WZUOA2uc84eHkFZEXIQv7YFs/tZM3oYynstmQ0OBiFBKdtjFiK1aDOHglmq
M3+fW9JlhjXqN+jUPcGe/MzH6x2kLzXRpCjJHoZd3nG9AUZ/t0nQ69o3SpipfqJp
S1cEIiOpAVDfO/HOHsZXWcHEqE+EMlo8IaMeC5BtHuAcBKV/u2ioc9krd3gbVqQv
NgGNQQm+I6zPvNxEHC1UM0cl8A80VLlmpYZjLGDeX+zj2WVyYz/CD/w6+J+0LLM4
BW9TpzrT/kM2LAAW3AcZs7uxdjol0siVQVXp6JaU3ND+C7I6UDzTnYu9g/W/Oo0L
XpyUeXBfOQ07/u4dwHAEDfltjId3/MZcIreCZelMLlOf70efvUYYAGEAgT8unOxg
5dlFJ/dEVhz0KSLeDUg+6Pg8/iDaSPZWNG3/IJTJ+Fwx8DWkUeKClH6yrtvNQ9sj
ZV6nkxJGNHXgG5pYN37uA+y85JXDkIgxMvbh0M6s8XLi71E0DGs+YEDX1kvERPhR
lIS/0rY5WAoCVXlvGK5pL55IyqLDOdjSWlx88VRnXhUZ/CpFZ0U7FX2PEBCqIJtU
faeWH3yRGaO8b6SdXy2tlLEtahCUjVEjDnyAuLM6MqGwWtCv0oDVL0Nl3iUdV4Di
Gu8gS3Kd54n3aAvTPTMSCrI/8kFDZRRGb+/u+nU6wRCiRXWBuXgGwsWFRhwjgEsH
PNxQq/PvBeLC8watpE6kjm2pHtZqLpO5Qub+FVwqG3MeRsdycwBEUeQVrfpfKcFB
+tuqQvhVPagGpCu9ls4fwaIH+u7XqUCx06cEmWB0WZ0+BLOUJH/WT40R7zeG8GtD
L+m2AvquqlQuCA+lQRvJLxdS0bi7iT6rgB3C/KmaZI4jyOnskbCB8R5b3+PBkbRC
jiXj5ROgTYkZrBbx3dsH+w3SrHfwKVZ6sp9jEwPzLoLVTcBSqh2mlU/5z5/nJBMS
oWK5+JKQ0YQ/UmUuwHzvXjV9NPqguWbkJNkHBxdoIk1jgNZO6q3cbzAnlRE35kxU
2gKjkzpM4wVWwnt/2COL57sI8jNY3lW0Ey+arzMhsbhb4NOkJ3LvuDAfig7gOh4B
aOLg5bqe/zVzEs+a7F/wxREO634Z2Y2uaaqK+dd5xDd02rkCSgTe30sNVesgUdhV
X1dVeOXZgZ+ZbTTKIfPwLEB7SX80DktgZVsOdFIkczfU4IWl608ADFRNVw4q61KE
GNpKQth2TZWw7gE6RNWH9fB7PVkdMVVQu2v3Pabq6KOA0IcfeQiYQb3XQMSS32K7
R285J+8NzdVqqM7uZlTIi0PesoW2DOEbdNuL1ffu1L3CTRJr52IE5R0VTeFX36x9
pwIPFo25yQOQ2L0//78Dg/tPt8zVrsKiD9wWd0TRWtqBcjU7tdfPmaEPK+P7VBtn
95+JZycbPnkD7QIF9mhqBrX6HB5QzzBcOpPvKBDNAEtXpQGuZLBK9QURl68v9CdP
Kw22Tfo9A4scIAol+yyhJVZ4rSc9YC43twCDLkj0V8iMIwJGtCAocoa5ebZJnEJ4
PovGtDfi95SRHRIhdWZ+JMYMj1Wv2VcQgTq0uEm3lngo04HlPUj3+13RTzeZ0/9k
ZE+PKBctcz5zjBtobZXYPsuhfsc57gTQMLQBaEKqWxy/Agq9xXmX+iJm1H5G563H
+5RHbSuWcE2qyfcR5aVuFcTFbLdLy7P3VNxapkBh90ZPl7rXUw4R8JLt4wGOhnzB
6/69mnUwQwgGUDLzF+WURZqY2f1kSzbOQjP1U0DdBVdvxKjoFjwVPeHmqHiOEV4B
LiGw6Iw82jiIWCFROLFLrdGbgt2wHfSyMQM23a9K6HRhDEgHBWDebb7DObPTdPAq
30PcVwUbKcGKRX7irjV/8TwoR7r4stUaadGH9fRhdaLq4d3/jVP7pqt3IkJh7ISj
5db1QJnQ4wOnBOjE8QV/0lAjXJoP8B2yQ/Jwpurd4J75olbmldhA3OuQbHjVfHGQ
hAiQT0nAk8/+jwGUtD+ywd4HeTpRp5tb51KElxtLssof7LUSwDB9MzNmhRlVfXIC
fdzaLvdk4Aa39Dj5stDuC79ttl+DgUMTAD1jQNG07HpPjsubGYnG/qDP0u0BIHwk
iQKmWvu578HoUYxa590EWEYVUy7ZTb3l9mByJiaQ8k8Hby3FO5y7k+FvxTcKDePu
+6KlQUmafK92Eg6BS4/ZA5yL+YsJHoz0r0l5C4DmjRiHsxOyDoBWfyfxW0aoYodw
/NgnoqJJNGp93Xt/TOH6G3Wzq41Ci5Ie7hvVNXiw0gpZTUUYLXwIinClsHnafzDg
WuAWjnc3DHlTZU8afFxOpZEzFsmzRs77Rt4Ka/RR0LfyHE7IecFZB0TyZGrqdEQs
aR0tHKuIN3hicgqwHmTBDKa9fO8Mc9d5Cy1CRnRFoqoY789fXVJ8UXISk+6HVR3h
+tZqU564leQwOWuxZj9eLy8y6babBpm1xNWKiSp9llHmGJNJYt1pwG+sxFnLaUEH
tPBTD3eKv/yzdZQ9lxfRu46i2o1IyKtSnlYNKu8uC8k+87MdU4gR8pMYBv7zB0xy
t9EQWoaBvvwRZcLO3CJUQR1BHHVff+kP/emsymSR6Z8RlMT+CytcffBeKDITPSht
RxHmDsEPnqQ8wwrIQHQX21vjxaOoijAa0W27psBjrmsteohOiAuiHFEiNyzn/jri
XMd/zLPA5EK+9wmaZTXBhx9AeH3dHdPW1VVAFMLB9haFK9uPfE1XzuIX6qtuj1yU
8PqV5nDFGpgJv1Vq2udratxjakDG+49dYqmRai2Nxd0Vkd/dwjWn5JOpjLRuY3ch
LntmjDTXNb00sqzCB74d3Msp3t+y6JVNsLyaNgqHqFDp816yfVEI5EYElW3YbR1A
fmeS1z1Xre2tTVazsro+K4/rWyjlOtmvtLREyTupUaGLNDcpFzG0ECASfdN6JTC5
+l3kkgFJnUtaYJb6SKVcumsovtxQunSNnOuHQrjt6ULVy+ma4FYSJfVE/gwPtpTj
Z7KT6f7gSdmy7qlQbLyBtLhATJuU5wAPJjQX0Q9X1aj26Sjunbfr7vahwxG6J6c8
Jzei3sAn5hJm5g6LMsAYIR2ATCoxJ4F58gYcqvJOV76lfwMaBJqtPGncdL1nA7uX
6afz7/YJG9r1Yud8VJLKsEw09z743gtHav+E1xUFJ1oYeLBKxWAqzEr7KBL+wsOD
mPW6z09g34rFX5v6Ow+iSVuYPIW7qwCh5YPBY/+K+YT6ivajK+0C7C5kiQNaP1ki
QqBk1UUywcOG48FgmLBlF7hE/tXaxPB3ya9yY7wNwGtD0dQoSfRcZaR770FGh8aB
mywP+DEv6Cn4RBClBeUYDQ0ACqUIEMkuryNqQocbhM+rXQP+SO0KoelbI+CFAdVR
XUteLS5t7L0p+6RxDGx/BkIn3RB3brG9/GxCOWCK6+jOWYeyZKIWBB2sJyt74E5M
giQM5SDLT7o68/sq61rE0VDLzsq1Nfglgi+9nB7NXsVpuH84ZY6eR6jtyjCl90rT
8pO5cBbriCqGMpGf9lN9POmHHZ95nKKvFgImICPXJaMqwXlt8a4b1YP5l1UG6/No
gNYBPzHwu4cI/p5DKudXvtTmhNqDFtY5lKMaePtzR326/szOx6hrTQlHVJeeF5tU
W9tajx5bKKnXI9JGHsP1NVLk2Uxk/Q0YMo9IOSabr7Z4CV+GB2xlwb3oZF/S622N
k+NwazUVkGrGWQmibEwnEqVJEyia6I+XZ75lBFxKE8b2+tk7twkHiquOUiBs4HQ6
cUvfEhf7BvlbdA6Vg7gypqELslHVQZwh5Es/folASTqZiidhdatC/Eq9fR8RiO31
XQQE3p30Pk3PfJkTfMNX3LsMUO14H+9MRc3hJLWcbfRJFRmOOl1e/Fa+mSsZ5T0l
UUrcLLEfvsmzsmLRU+OMqkGHdLtFsu0F1A1yJJLcFRv7YZdAofaJW1pBGOG1rtLz
RUyguox9OdJ+4eUJkmBICG70Er2uHaqGF/C0qYQ9361h1mnbsg0VjTFE1h/V8E8r
sQvEETglBXWVBphpwp0fm+kel4WGH69+e987A6cEJHvJgZUTvdq1TGbC1LGzDm4D
7NzB6eYuLFCavGRruc3DC5d6lqNo8kVV82PE7RcxQ+NscMze22jVYS215EStCLDo
gvMFT2LNZOsGacOKLpav8k+X7rtHNKOF3qRw86ye4h7HtZscS0r/r/wRzEiUlGzS
9J3xyO62Mr801tgmBloDWmnS5Ugum7GOXsnSIOeaVSnORC/iavpiXsIwpkiZwAkD
pPCs2qtuPgByN6jaYp0yWdfIUqkGdLyf3G1HqnFvOZu026pZLaz0TVyV7e3Ir1/u
4KFWA1EcPtipaO+p2Exoyv84Rch6NRfMFc1y/GI6fqKNwRDOMmkClRwgrJY34Gzk
vxKNYEsIEnFDdt8WIGoa5CBLrgwWw5ZDju8s+thE+ugeh6BjWXlErQyjXKOt7eWs
r7tjVKzZ9d176jMnNzmy7LJKcWdoSyMmSp1IR3WzU2efsOWjsCFG8/mIqLhm2Hji
6JdvapLstXmdkOka6mmOsKtupWd0BHfypENhl3GV2uACT1xuLMUb+ZlJfodsTPd1
hbIj0q7Pyk/iKrxdWaHAkl8uak3jfrtoORHSIlu9jymGd5btCqEq6i8CI0EypGH/
haLolzDP3ieE/tfCQQICqUwatykjGCxUlCPCOwnLyLio2vk++YKLnSsSVnRE3GHk
t2ALvLHXPDNlhpt+FobvmfT5It85y2WwsaljKe4C3aMoqFLZvalN5pZsWolbRqzM
Xpuu5pGYm8tdNJSgp9zHB2QstgPTEAYyv1dX4w59VHig+b9OLM8vFS5o+XW/iyt4
NT+RE2nVWg3hqM11eX4khZj9EA3YKFiyGaonD3hC3jY+4Vq8BukzzM4bQ0wdPqE+
/43llRt1dGeZKHqaNdJJOnFazfTb6hBYcNotLvAJS0l6QKBNVAYJXwX2leeA561f
Hocy7ijjnJ7AEHLx45LOJLIuhkovlIsKPxway4OEWEuqyzlEstuM8efxqkTdc7an
p9WVoK5JoP9c0c1esgk+rj0ZFwHk68dcjXOx3HrdpqK84Xz4+Tkp6rWz9cxtkbg6
9VO/5srx8GouSt+3S1IAnmbMHIh3m+fEMFfXeRqS1PKtwcVh0xTcfmqB3Vw4B1e9
1MNKP1lCKCwDIXo1ondumGZYT30W0VQ1bVbZRB/5AiPVUSqxnV071KX5akmeNa+u
f6/ePATvjNjvltXp7upGLsW1tRR7GRKIEdFUhbgMrdoaKkvOH0irJBsbEcSMdtKK
IgB36HXr8aJ1yug3Ugg88T3QjwCm5tNcfSYy3lYiuwqfRG31oclpYwWAqeNbzwt9
mrUXani2d+dyLzqXScvSYQmbSuOBM//io8gYngVRBZR0fp1RxKGmH4KksSIAf6UO
jVkI7S5jSNeSYWJ4ywpf6cASWTUK8D/E1gCC7bm3KiFNSDrznsL+cP9b5zw9GPHc
I5+wbIYwKYXtGtbaKoPa29m8Sukwu3J53U38DHs+PuuN3jhY4/hgRh0+wJOw8geb
gNz32lsZP3XeTH2F4tdw6EWbX2gfbEC2y2Y06Ot6wyswRpnPY0MC0gp+N+iZZ14J
13N1eR5HVfnLsu8Hlg64FE1HfVXoNdWH7UWhCIjCuW0Qimqzqg5utEbeQ0HU1Qub
Wrrf01JuI8o3+9ZStG2/bSEabLWrk4SyuCeMVpwKz8TeZHXyPOIIgv2jh0UfCcBM
cVc9a6bZEA2UOMekUJu2PpHMAcFJyXPRPEvsrImmciEazbF7pynDONQAAYIRRtqA
wSac+dOu+QEL4SVnfVEheD8Y5QucZrAwe1MwmQG8Oow/XRyncID7EyoxjDPDIwWa
1zO7mWBUmAoiEfKdwx6ZbE1fa2EEjBmISQJjG2UXBY8yvZOWY12GiHTS/kJTtg02
Bzc8G94wQhuf8FgREyucih3BekI6PRHCvsqMVy8bFmCNvkDfxdMmDG9Gy8fcpHtx
izmjAFqiz81CFetrfuFgE+fGyHl2A0Mat+dx/pYO72eB+3fEmRjR/Gx6A8bKqzeV
8ZBGCYAr50UkyKzILCt4IT0aFVQP6AQali0HZv5zrhCMJEs1M20VwUKo4OBbUdOI
+eIF/HlbvdutgWwFTlNkWhWwlLENAUzP6mkvXPBWdluhWJIeUrs7TMiEo48UsUUS
F/b+ZUv+YAMiMBSpRaMKtP4Ikv0EhqelNk89H50NBElAGAnb3wneOqch32zWjufC
kiaVdvYEenQ3sn5LDs8l6Z2BRQEa85yOhjPvrGoZNTI0EN92PpAxvtxhm/ZI2l6n
+78BQZDZphoE4JYpfz45Gk2VruRe5VGfqhsp2/3cqINieajClPJLRFTMjzAySZQ1
Sq1wrARjlw6klNBpcxIBJk3FjFnO+6qA5OTbQ5ricrBTpNrRVMZE1URByO05eacR
iSC6hnNyJWRFsIiPlW4bre7sbOblI7e3GhegMvXiTX6KEdyWTcF/FSM4kG9R4rnr
aXQLS1GAeGH9WX4dYzYLtho5XxQvRXwAvuQujL+JAbG9pBOIOvHeEbe9FSrzkuvp
9ysL3dGX6OUNBXsJnjyJFRUkmZJ/4G2d40g8gZ6VvSm6CEKbUdZjdtKVuYag2s8y
GiPy3rtuvgT7bBM+nHJ4AjotO8azdlxuAOHyGFYVkENa/ARxJ5Hvh9DDeslUmCGY
l71U6HDn1C0TH3TWbV3PuUBzHt+oNTGNuav0ebF8kPuB0NkNRKbhuMnf+xgkNBNK
c4oQYtXH4IMTwL4hAnsHJEybTJzZSQTq6etnaNbY54AF1C3CEe2nH4QQl1lmjZNy
p41Gz96NxxlmUAy9FuhZxQXeFfVDTAtIfXVt0T3zA/lJQIbj3q1nPvpOl5itNDpL
Euku9YkVIOTfcXDfOCDMrHh5Fvo9LVSCiSZuJGf20XHJbFXzJIkCTffwkESBG74e
RWjFEI4/WAuk0mT3WgFmj+CmtPz3n5/c/aaL9VDUINO+pIdlpl/QnwRKziSUd4NJ
dMo+vXWmHjwngwZmGBWamJ1bXAj4BDs+S89VWLqplk+S0Opgdz2+swviV3o3Oz3X
mxyCHK6mniUkMGtJVtUYphq7H3PLGswtcKTd9E+/aXgCrjendahbgMpnwb9RXo7x
Jm59871zU6RIAdO4ghIo7O02zTWZfE81mKgxUa4j4Q3xC0vQO3E1NQS8S0M0VSdO
71Mc/ZgnACbxB2j0YCEIUxpUX9f7JrlNX9Mx+eQ6/k9VEVVyqjvrr9pPPMResQRb
7EHDMPVaPkydW0mnIaWyzojaSW7IhO48/tcfAdCBXhYUv7ZhM4hNXXjCngERU2f0
bD+5qonPrUXC8bGYlCfJ2l7+VSfEPCwpJRQbl1fODLFejClCaOdk4iq8aLgQI1Ct
1mYNsi83ZxUL5U0YOKb0J3OimTWRqSVNWWA/YWoTHNHkHwQy73mUhdP7FzkBKu00
Ne93a9k8QytJNSIs/SEiFh/medIfmFkjgwtOUZSND0I+czuqXb8/oMvs4cfInG3F
acy0X43fNdqwsxVeuPHWy6slTOMe2z/r5FdJvmZtxHzXOT3is2eat4WfVNvsWUn/
9IksxC+H46wN+sZJiEDNwd0lRMr3Ch4v56EgPkvn1YmSNL/rFStJ0uxIjviq05IS
CjRbb6xygN1rU6xc1sMIorKEZi/6RXHGlu6ltDvdjgSWXhIQ5RuYupo7Ek/GJGZ1
C45tfK/aIfjZadil62m0AI5XKQwlFWDXfY8rexE9ltX5UFT58NbDfmrp9VCMkBLp
t7ZplL5APJi1XKhnb0e9UgXh03AxN5XgCo2ToB+0ltW2Xw2OxQK1C/TJdIsumlt4
omk0rBOzI+DDwim1Mw0sfZYa2CFzBjziSLvM18MjYY6Eip+jvsJLeMvmy9plIFLU
NqlX4AHTzzxyKfEjGJ6jRLym/Ya5+dcQZDPaTO8JcZmwt8E3rm9LbFNFqjNEyg8v
mkvMP7GkRM8/2+oQAFwAwj/jdUNOTi12a+Fm/iInFDwAByPao0uuUntI/my1g7bO
u0HvYYl9M8iey6sb5trZBEE5hZ9UXGZcUXFF3RflgdMD7TrPbNT2aoW9hUHdQPO0
6eKxT+JIh0t9Wn+CJV5iYsJtfHHmICSxRUr7mtQP4qUrFuLllQr1wcEQ419W7Cd2
EtQrWHYkVFM+w56yFnlPdhWxxj0bxY9KgHRrFCtVqA/37FqnXx3LRKnKLahJc2Ul
iL0cSlf0SXwEzwknUCuVbuUj96MLwpoJ0LCvzmvqKiYB7VZvPAgJYlyFvyqK+h9S
WVyrYr+lfCLROwuYqkBtaR+HV3tcTw+mcgl5jN5Z/n3SZhjNcWf7V33KfWmlGuEg
8bDOHZfWcKRdFsJOe/iJXgDqV4yh+tY6IbcyR2O3PsmCMFNJELCfvGbccjBKEQ2F
DlOCh8adfwBSQMoAHJdNYzZUGUZAGHgY59qcc+xozoANTiyuhO3Ez2u7/ET1NjZ6
jY8jGAlZ7fZvdoQMpV1SfR5dVN5iLrNUQ08hgtJhETm4jbrvsk4qROdGVO+7LCKu
c1b4z4SBqZAKqC33aRZBXerqe4+7YAUHyhEa0s0GHyPrqYTJr6p/ERfvt8mcD3OC
K4GSSMr6kaPHgyoKEaPqjt9mdt5RefqDDz+XKwfLKGyl+VDfS2/heua6BsUrCHOp
/Pv8EUsZpulUd58NLNfXf5eoeThRx6SlScv0PAs4xgBQce9S0AXotgd+w5xMP1Id
li5pr+imcafqp0hNSi8SB1Lus2DGcc3PvYC3C/zg8/p7r6OgNw9Ua3ZQ3pGheQpG
FX+2AjQ5V3/zfNXCPt6XkDN7MY0n7mwX/jjO6nXmND5wAew1LDSDmER/YnROlarS
K9IVaaVV1aSPp0UxIVbCg1ykShOw3Tx8J6KB6G+cpn0iVUcw4zmhb48eFrvhBJGR
Vj7irZhHf5ni5DELIhoCtGmcnJjPsuqjHQVkpNC0qnRv5msaOZzLAIgZGL2Nq9hl
5hzvC9ztPgvi5dXWEUmaAxea6wZwg6DOIdJuhrd9vyzB/uuYXEcPDyNcz196ZgmC
8/Dm1R8BrkbPv8lpfZloKXj6LIQ5H0emWJAxOpdPAJNYyCCOC0J4t25aIoZnVKnf
sDf2ZSwGFIcPQMuNTle8l8ghkV8ISAYvLU9WgV7tDRlvh6BrnGa8ou9fyvNsvHf8
qMWrNDzR4UaxroPe+yFUG9494WONnHM9aN+51VvONn7c4K2imkGWE4UIQm+IeFgz
VR8GQLfER1y9AyFktgyHvhBfFkqZmqa8tfIV3WBHqaDOVjsMbsmfl8ZtOnoT8QNI
1E43aWVV4b3c/mKR1b0tAFe7kJWCeYRaVZp7eWtkRLgzZW/wmSNNOyy5Ov6JjFYL
qQMvekOh3fF9G55lCtLudzHEzIJ3w89cF1B2y105hKw5nG4WlnKpFICsMzWVaKWF
4oO3TtD3IP0lAKBSnAOQUt+nbGlNJnGZ3yzrQKk6GZnyNdQO0EvmqxlSt5qsLPIH
2FFUz8CRkIHTfS5qLVEG+TrY8jKP9/nU/YJqYTKKxFK/d4sRca0oBFpgQfcFG2cV
kYo9YC1w8viC62D2FPSsEsuTlr4Qjjths36P7MKJZ1oKsCsGWnZT0Ypn5LOmp8o2
VBR6WASFtLL0eyxugHfVjxBCtdkhFO+tzi3eek035Zh4maDIaDXE13HpvM9lfVVo
YstklKBjPggeqywhnLeKm4G5nzZ6S14AEWgJFDsf99mv9P0blcyhUyAidQF/RU4A
sQCQL3FDYkFAJDiRrNvj1h8dys/F+U7PbewxxXNAFj7ItAdSpXjFfxisMQMkFIDK
tFc3sFttk4ctdFUxloVodJjcKYf4ufpxrAMOyWi6lX0miZYowmhG0CXbEGAS5aZt
+4997z94YH0FMFy/NdgxbwaBFpDGVPrjYcOTeujk4JA4N/NeV0RE9Nh+jPJ+sMck
8Zythbih6y7WHv95Xr/XePCY185ib0T1/jzsGcaURD1CTgrXrxZQjpHgpo6a1p2X
xi6bjC0LWpAX2aT6FjWcscH2JxCREXMqkrlbMmGTMOTKM8DlesW0kwXXUvbkBh2z
JTPUQcHO8zjX/0KdKbdaLTdWK5bGvUrlp39RVxUuJ/JBlJMnx2O0LLInwaSlQI8d
eBZ+2BASsDs8594AaORkXyN7XFG73yhFzpvMmm3g6suqKZ1WvX3mwHpfX1DPjO5+
8rzZtdr1JaCYmVLVwkR/AnA0fYXAm7Y5hSe00ewEXkCHBZgsOl5U+uQ4w60tq8M0
xvVUcEG/CG7e3DNf6Ytx3FoqOW7+2AC3qJJXIFWiLzS9MK79B8pM0BAF6fHnEo28
hRJ5xnbLil+y69NIpJFvI39LHAvVFDC7CIuqNH6JJ6m9Yale+72gag5qFmmxPe71
MrbZK4lJom55zXfPWcCcDGun0vqa64mZPP+aaH697YaHg2RABmjRJhk3F/0449yx
tW9Z3hCpf+f3+jbq1wM5Ve/NqIx3v25cfQ6KM7qoqg2GZ4qVmuBMHhvr6MTlpFHb
sM7K+NxD0iWUCAmf0qScbKES9Wvx6bumL56fMz0rDJ2SQtQQYstJN2eHOFqUo9oM
E/vIFp1nwy7rPhRAFq/vP2tienYpG77PDUQdnETzCvUWlhpwPVLOQUbvuHUqm6C9
jNsfv8WjdGM1mHd8ggh4QL7/qKtAK9vaNeXVL2p/d6/MzhyDp97q3V2kXhJwnMlG
IjoxQooBTtm8dPIM3qoCA89RyI6wwh2De1osKRyshEA7e7ny3zi4fiP8q6v7M9qC
gGpAwnGAQ4qV22Hwj/3dskd2j/H6zbMFrEkASOpRUPb630OLnWVl1F17V1TEEGiS
cXbK32lq6w2gIxRWfMKWMFQYh7moNVZibczuGC+JOb9uB2oaYchJDo8u6v8cgGJs
JZ3glVFmGRJnivDALzv/3FqGTpChTbJkQ9FWPug3JkigZ04vtQPFTZaJy7lehjGH
EqHjpn0O3psSrhFVk+mlCm9H+CZEMcpQv23fzDacz/ELtR1zKzFoiguVjWI0fqHE
Mn6Hqpc2JzyJyZtRYmnHB2nmP1cFZDwE3rVU3e5Ojag/Sb+VxVBBEXXnKP3GI9VE
/E7D3zEiGzJL6c4VEzhXmOnMUMTOu1sC8eouVXU05e13XRju1iBFasaoLRQJm+fT
O6j2dcFTDs0puLdPhX13OLfeP7nN8NmA/tlTRJ3fnjA7yHsmtDQy/v40CB1fz7KM
KpziNU+9qefDmgxMy26jWujyQy02c0F9lm9652E4ec4h/jQN/paS12GWJlg/MorR
3yNP044bH1gAC/FX6YtxeA47fTcpBW/ZGvyxuNviTy81/AY9PPq2MX+e/uhCedLu
+622V5e68mcbQVAM2KWBtjuU00LqmgHDxcGvUvf8lR+TPp1jd549fTmgY3ffx8Se
+xrLyjmGmwraXV5T/Lr0BH8odlEop6gS0zFJ0cOJibkaoP6MAuLOxhanFVa2r46V
Kufjy1oLwDPnkb+MzMBePt8XizrLJnNmYlj7Qc3+eQgNfxbreGF5PqSa8r1AQpAS
73RIDxNtIWg/k+rodOtBCh9B8lW1HkuCo8dbo8tLOE83A+aAaY0GPnlwL0jaoPvr
uhEB3maOm/cq+Gb4zrNX13c25t+nLBoR7IkplgPXMioy4p4E9BGc0XpiLzgSMSkG
5rm6afl7cmZIJmxIZbrxSLq0T8dF7Tal/er3mCWyXK7zhjRHIIXBA27rTeLEFLnn
9hKBqG0WRbiaGp856E/2hxqFRuXlN7jf1ykahkQIY2ThYODs3dKD/ZD9aw3DDoSW
X9i1kuECsq3wbMp9wlA1WU1+yFwT2EKpGN7SdjyFYaqXz50b8AkIwEpAFcUhUV3c
Hy5hWpY9pIsxAm+k5xCx6KmeZxlLioa+nDvWAk15k7eR+oTcJWq/xHwhnt1l9MJF
V8tAWd23eRwpCPQvcsRYacbQWVwa8mnhj17BkpvekRI+DAUAA+zpSWItpgz0bWiP
9XhgPviHN+nXgzIE7+UOQjaeBoneANq8ooGnML2nyeu5MVrSCpg0QPeFiKAlFm2W
eGzfzPtzhTfwC0e1+ng/9QVbC7YR3Fa2evGZ6MIe0s4ZAuBcfG2sKZ39N7Ro6wjj
Qi/OS0aT9ks7A7JrBH4Fjf6hwZgY4XDNNInN8tcy/tMwLGG4hRZAt9ueFClv91W7
s84+nlMVu0v/RIVFJlrdX2hHmFaoIBTKHtfsLgSN/X1th9p0MyK5Xn2CvA/I9Tzg
ceuTtb97Ju2Myo4tGMYJPz6vlYO4Kndt+cIB49l+L5k/JSW5f7gqKFm1y4chNDFm
vDS2QL4Vc1Tg1MgDA07/sQWp6Kt2EygsB6AB+N4PrUGlEoKS8yzDsbnbq9rt+f5p
arA4AsOfAN8MESXw/5ydxRq2efRcZyydsF/BM5pKYY2ggJfCA37VA2KEKjzw2Hu+
RRkht/WN4vlHjrO0KXJ/5uU3mNCdUOhpayfmTkXOQGLvoI0IJ38iycfBAztNR+x/
R9swjCOluXC2snBQDIwMnc4pxzFuLx8/OoVO8eXQIkz6vDLfkIEdMSuhgIKb40E0
kW3SMocAEcipTzp1Utf93NnqahQL8OixsO1yBu+CcO86r1O6IDyhzjg0MoXH7MQ7
tbqaDdquUs6eeOFA2BbLOvwntXprmct2+pb8AKEe2rz8bEboY+FnBRiVL4IZEHLC
xmR6PkXygGUCE+uKWfZKLTQcRB4o9k7nvL/qNRBNzl1/k8naNghRLQeekJkZRXRj
jMIIKzIvjl5e9pZfnch7W3X/FK1a5Y36edCrGkRD24cI0zmpLhU/hdabux8CzdNB
y0VXHOalkx7g1XrmxEp+2UkjMFyosDPXM5nQGkmMaFpLWa5ELPYIg2+HDvkmaEiO
4FtgefH07GVsgC4w+pkd396fNut+Oz4yNaJR4EnBlJqGZNW53j1NU52ByTLIRvRb
V1/PA8luZhsAN1JtwNd/P5S1KSKp4QkYD7C+jkqrakRp1BaapdKylgeMWQcIOBPI
/WFGULk/TlJ+wFYq65Uh7Uq0QJOOMMqcakm16eBvI/ahGcW9QLuQg6lRFNPtnH3m
5R60LeaDJwXEqZR8eQK60xr0bBJsd7x3R/3BitdA7415JaJDxv0xmGf7pLXSX3Ew
aZD8VGirKV9Y/pm+oU96nCSPrOFYKoKqfg7B8OsyLWrGobSfrQyjuHhlm2POzcE5
Zcwuvkt2RHfzBsa7xAjhOh+hRn27QRopZu3lTgO6oDgybJ5+Ps/YC1Gb1NWfa+RS
RnYEgKp2DnML4HfiQfaelH5d9ohqLGfv7UmF0FRFioFm56wXg/0m/8GfT6JygeEV
x7vlf2lKktNBx87WCxJBT1uXVpAIF5lKytJAWfN14mFpFpWoDr9QlqPlIQo30f63
KmvzvoiGhZhfKVKiu1VBryz40H3pUhGyeNhMo0GGRQzdK7Q9P/6ibhRo1LkUHPYl
rqivZ+q3bA28c8mmIVToiKO8eYtDnFPo3lWXw/LvIlL2lNtdBvYilbYsErFOOToK
SjUE+iLxqNLpVXvKVy7hn37u8HIVI56HGTe6YQ1gVLlHUE3lPXrD5/ALaQ5P1vzL
ySpornh+E1t0x8KwKI3fzzVPcpIYM8ocuLRQmJRzfhl1YsO6DImlBwhAC+sfiIyO
MqWnKb5TUfyWWU9uYK+iyfhUCtnJqM6eZwbaOe9+Z9M5FLEHSVZuGJt2srbR7m2j
6pw6zQu1P8zHWtVk/1tNdcPksIhEhCQtQrJ3UIrmRDW4A+xf9fXxoKJMKFRXPFOo
0ZEYLubPR27gc2Ln7u00YRlTsOtdKkUASwx+k6sPV9+qr7G6OLN3D08PGxpsH2SG
Uw2h8T9mCYj0OCeRKmCvyFTZDW1j0c6rkIxugAAJKctHSbJFGz5LR8vavGorxW09
p97ZW5Gftb6IOBe5c6f5aXkU/rrbYhX9PPPVYhc8R7njdGHqsekXoCV/Q1oz1cQ4
J7b29cxebaW6Vumc9rRDvdN40PANjzeaYtKXl/N7u5Ajj7lsIsGLFz15e6JZCMts
1jWe2EEgC1lsN5vu7oBfMEI6Z7PmGSI9cxflZKQrMDRrAv/IJHYA5ZIpk5EpMoWp
fr0bdyzElCbKM/7k6vd9nSDh9Q/NKtFfBV2lud3vCZD4pVMTORyoAq1f5LQEYdzT
vyi4A2oNXiv1BpVUzmDte+zUmILWIc1++PerJ5kfyVopXbZSniWd4MdDaytAv9wN
i/1KGXhfXocGJ86I1ZKxU7rKUEnIe0iTbZq+GqHWDRu94HT0y30d+itwFIMbcaYR
ptoHZtGN3aqXk7Hhmg3374+T+BnvXI5YZK/tE0j3Vjr3dr2j+CGsG6GqhB8wpPz0
8eZ8DDRJog/n5dhamm/h7jWd5ut9g6AXxRR3FKHCuEA4IzcnN3a53PCoPGf2OrID
r3HdbG0YLVaZLs5OoslQ1zpepubnaausmAsMY+EhM22iYpYUYflnkuXJdHrRgnYI
4x14oC3QjGdO0r/uqrC2bMmmnE0wQoU5oWel2Lp2DNx+jMkL1oDbHG4XMqLUAnjt
laXvFG3JTlowRaySTUZzmdDsnUB+5HRWVKxEd2TS/04TM/HqZxkYAFAtsk6fl9Kl
upDWLyVdgbmZzjZinH+a75jBf/YuncQM41pCQGJ+kZxXV3/450zKxRT4idEmMYZV
258TElFGdpIeGPWvSozNMfgJXupnWzxbl8oM1jgILnu78Qf6b2dP9qK5ZoR9PnpH
DKTTj8ieJ84gfK2S97tvbviPTsNnFPuyilnzaDeBzmAyBpgy1ZBHfKa73M92Fslb
BlMtehpCqjsd+ZuOM8TF+wZg0GAY4zQFl+u3u3ABzvP2eytRmZizbIENgsQaecfz
TCkGy9xXFFyS7YM0N73IYTv2LZ05wP9WZA+UdDh36gDdd/trLTPhsz5vXltN42T8
XD0NYhCjdVzDon/lyOuJwlx/HJIlZA08P7o1gOIqTt64N9znIL03H04pEBlGSl3T
UqAbi/9G1Mf8Gq5sYwBX9S74yruOTZM3siH27yCFbed/Xl5sKRNVeQgKRC8cq5AQ
2Tbsw5i6KUNYNHEgYgitop+Ro67HMZ96WES5m8sXJ4SRGi0wXYrI57uzyuG4WBMX
zQyGbgrxAANYRaUh+K8uU7gi6j+u3unzbuwV372rS/to/jxVHI56nccB9j/Mh10o
Xx5Vmmx0+f4nfFsc2Kr7T1+2yiXsDhSdRGB34IIyVGLaNygM3B1yOFjn26uA29xj
ZKmsbC/uViiGMpqAyeQ5JeTWS3BqpkuAUm+GQAHCXcfhryypaoXXs8v03orzD3nz
fsXOqi/ZHF6kHpbNt8/CB5eZlcUQHqd1CYoHMLJDSoOGxmto8J89C+FkcKg1YP21
A1rGwyXmgRni8GPy0KDgT7pWWwnGkrvIf8YIo4/FQqb/7T99Pl4yVKx8mEL+OGkn
SmaJ6kvjkwwgVcKsSAgYJ4FrdXk90JhBpZze2DjAfLfAEJTEIFGH5gNJx3t4M/wn
RBS/xvaia6hG8Ia0YVwIY/19j9S7RNWGrh9dnxvnNKKGAIV+Xi5AOCs0njOd+MRO
qOn3I8aVV3ye+fIUOLfZgIA3zqfRTdm9ZtEiZfqBqtWGATxSncUsIbe5l9hCybxh
XmXJ4LzwEcHb+8UlyO6hRIvs0PGFtVOdQ+h3QY/+1aViWgkTZhuMms+LCYmqFGlW
1cjJZEi0mfMTQ29WojgsRzKdlAXNO0CZN3/lpH3e4qdnvUDXU2vxyA9q6Yt7HmGf
dVYaaIKFESXjN8xe4wYoQ83wLbgo9lV9MspVMJmgucUd/tHQsAOre+zR6RZ9EhG5
HNpNRF67BWDkX/lMmhZtWQbxSMPdiK9nBArx2hRV2tG8MxkWbB1mbkS+5iq6cH7B
FFACXS6GtcAfjV/S9qRFzl5Wg8usj81zydRYuaCZEnnvuobvpUqd1ThjYiN2qQv3
NAr3t5ZxEgjXbfpmsIls6Xui0DGfznF/HL7TvGJGqQy3M8FMe7+be7etkFmQ7DF7
yMIPj6XTKM79zCXsUBB61O9BtuQU/H9pWvlNgnbVfcV8lg4X4dH16xwuQJM6XBoy
Tp5P6abYgkiVBE1H0I6SBFQ0yWL0cyyzGH3dPssyVwhYoHeKouRaUZjOwdIIeXwD
Ht2RgOYVsP7iFyrsvPCQVwX3dMbZ47Z3okPCfxWdvzmhCFIL1DSGubQ9Yyh+QxBc
s2Nempq0Sa7TbOYbv8AUkkGDZ7QCen4Nv8wWIm3Xw8Z4obRCQZ2K8kxKRLFcAcF5
8I6fOTIrxS3hThFbew3wr14YVlUhIKvjup0AJIR+xnlobyh8FGZ1miRnk0z2dozx
+jSkQSzDmE8UtEVBIT03nfcCPyCDVEKsiVdWvzTHduUUCVXLZVg9PVMka9pWPolU
I71ESX8kK176C+V4Q2VvK9m7lF5/bIlmtoQoPJe6GCuVpK39gqUBvkcfrxDqKI66
LidqMPY09geGKIOPRmLHVjuXa/XnDnXBQSYbWunePIhpj3SVE5KdJWo2pFRhhRIO
9Pb7CfUe3T3OyA1E7hheJeTe+OlsLdg/oh1mFN4Bd5YaamfHPi/WSFWpnMG1A8oC
e4dLWRutcOQgKMLIFwoUu2M4mw/qrd6wwDF3oh89eEK6t2EDfQBqfNlUJWVfPtcx
WpCqKH2UbS5H+RltAPx1pUAHfqXxP5nQSDZNK+FlcGKUxyEQHnCD/LzhVB5a8RcE
wU0w10XIxCpUVnNw+ekUvuuU0NxmNpoNxrp3SKPDDNBqThphqiNDgX2l4mILuv18
yddRBAW9/PMmRmUM9wN3jHxHW+VbTvuLLsFqK74ic4admloGSLd65+a2bPfZrSHF
8Kq/r22I+iyDM1xSsFHvWBwFIvNHrt3y3twZgkgxzp+Wo4xJH/nrkxwEG/4a3iSp
HYVYjQ0ML3Sdm7vbb7W0L09aiwYTfwpZ1YMWjBEHEbTobLHkG36D7Fj+F/e0ZUL1
d70lZYaArRkLzm0GkeDeia7nRgkPpxlBNCdzugRElzMtey0rKJqOP0cahdDNE7gs
RI0/EOMkb6djARV1o7StfxZotw06T7vRZouE1K4pG2pLJ2j+0hnxg6SjuigmlCXE
l4718VuLNZuLsr17RvfpOp8tSM/Ar/EGDOyBGf/n1H6x6qQPaJZ7mkBkCrtN3twO
RIZTGKTnwDpstulr9USBDIaNha+fyFq4ZB06Pgk24omMMLXc7/3bn13MhwfX+1Oi
kboxfpoumQt7NjllEC7r+9gcNh48H5L+S8BmrQdjvEySU31M8rFWLecYT0VzXY/X
Yfu58GKKKwFTWc4K4Sd+D57SMISZK0l7q39PaQWB7d3OOnQv23QOf47upAszRTw/
HUX+0UMwimcJN55ITrsMQDkT8DsFR2t91GPoYBTlDv8wsKxmQ+frxoSt2r4wQQND
cDJYTDEsvpwv7TcdNp7FSyem/2KnVWezLYR03dDC8raxKpcdnDk2wSrYniEzLiIn
oOezSqSI67iq000rVjVLJYT2kCuzJt0um/oRakNH7fggxz3PFZGOOtNGEnxQm91l
xm5MV7EhxoPYeA7szho9fhIwPkWHjyRNdU/1e3qcl/ep7mY6/cFOidQLs5GHz7dw
Uqi/XGHOy9EAEuogbD8S/ijoi88trt5uBFeStdid6MGOTQvTXpbLCdMC8FxNvTtK
uoCXqfXuhSvscvbIZaIK0dCgXHutRNKOBOmUQbpOxYG61AsSj040LkrClK446ADW
TQs7Zrq6aNPIZOCejL9b+tx9G85JVZgwB8V04yaT4p/s1RVSj/34IVrrei4E6RO2
cDyKHrppJbJ2oHPkR3QRt4EIWvfrIkqjCzdYVp6117ctx+yXNlfwjN0YhV/CjT9R
ddb+4eOMgIXUYM00mArTu4WO6ffmtrIXqdnrbyieXtsTNEEieP8ou0YeZ6a+RsWC
muG9NMjEZipgzODkzaUyTxsi5eUPXZ8St/q1bP5VsQaRVYhHoQE7pl7SCreKtI/D
4E4U+6w/o22T04pYw+gg4hptUl2D4xY/2aVEuq4CwqhhavZrYXpcqvjjBEODW1Uy
cw4Gza7OHMYxDQZzsANkxWNgqAzlEmfaXot88IgTWHcf5VMD9VJdpY6gRWujMU4R
JX6sdZBoAFnXg4VzUET2gFdyXP/ca6m9gxD49Ppx7CCdHJurV+hPrm+KPTo20zZ0
V/mfDMeM9efvlFHeirW/X6FpU4eoiG+U08zo0DqYUyBZTrgFXD3L1cclfvfrR+VH
V6il07lL1Gc2przCgSmJ6uZTydKbGwNrzVpXPe9uc4NjPy6KKUnZ4WjbcgxqRr/v
+a8EtaOuFEXX5QEM3szT12l3dStFDIlU1NV7OATuvzJBxVUY1RESv893GH0o9qA+
xPDcLSct+4FsJKIa27s8+CljFPNf9eu5a+Wr3IyrsMYQcEhMkCkQCtR2uY3x5r7h
R3YkFiYd+k9oy3hLQZ5EKkFGL1uIPLPX1BanI5MkSOYjDPkzm8U0e9niFq9+kKLF
tU66EGBAjGWycqktxD8R4a6w8PbKKYyZvaeM6C23/SK0Cj4dkU7cN8t9zzbSFF4U
+0jPv2x/dbXfZeQg9+SImX40tZDIkG6rn8sDHajgeOlsNZF+ooiOTyirXDQJLFn6
35a1QjpNjQijfLHbIvvfrbDtI4njdBFgfV/kASOQkN4HNOAxjTrlsvGQSDQT7Mj5
vjM4W3Nqa2F4r05xGgVemjoJDziAs7QdaktFZ6f5qS/mLmq/oGqxQSCIwQ+Cqvua
9gZ4WtT+9eNgxS0cSHtMerU36nLnUC7XeH/9TLmiw948YQqhkRd5bnskOmVHlY4o
LI23ig7gJXe0bLlvPFdPDGsOsQ5gBxOq0UISZ2hdHQaRsQwwemT2mrjg6ausx1G8
ZxXB04SPKPGHLcGRThHTCC3BzX99O42YMOMT7y1LqkLTTf915B+sL9fQ4jnQvZsj
Qm7YTt18fUXbeqTJFUOzm1ZEoWY5sd5lRnUxZgkW5ZHanDgfctarcyVQbA752uUv
vR57v0KmUl0Ij3TpHD17CJ3ZUGunp3klU4hoKtZNpcPStOl6xO8wwEMf6X5srqY6
MOxT9biA6avZ83aTyCu9SAgYZ92gNIEvKxqb3ODGWm0A0asu6kWmQ42VVekpXzqA
D0fHkY50Esf0cL/3d/48KT6V4bkdvhvLuO5b0g7gEIR8X9CLhR1aQNWo6tby3Cnk
DCk7tVvUONnZwUEibMeZ5288SRR6bDwUeHftn69QYmRFkFfTpRntSVEg5m1vWO1d
4Y+5GKg7p+g9JKbEyYV30rhLj/BOxYaD6E7YSSq42Y0Hgs0XvMJ+SD/EudT3Pnw8
jedKDpudLPnRkkG3G2iAXGYfQmnZfPEZhnpJwd4ro5WSz4G8XsEhk4kUO4UJKuPc
Ncx+QVXp4m4lEddsbuo1IM+FVSq1tR2FHV5uhfilOEx91fMW1QZTCpJNZdWL2DZJ
bKNhMESQ6tK+sq93ATS9wMkbID44DSdG8VYpuZB2lCyO4Wj+AgI5g1+NPZKdgc9I
EaibJQu7Eec3aemou4Pmx5Ci983pUKgzCYTLcrAooP7VkxAIR8vuf6MNZeVQntrR
wCX9b4cEHiVnZMt174wns3sgAT2JV9EockT727kv16lLTqwW+3YZ934heCi6hBex
80FzAJq8i8w1mIO48bsD5QocQn5Yfrn10mO32JUH/2LHmSal7ax4vNfHsOYAAIjr
NGb2QeloBAsM959yuoY0C4CAs0uVf9/Mqu1lBQwFcLENpNoWr8TbnFeOnFJtw1Bc
V4YljwVVtqK97GagFe6VCvAc90x0xAGbuQrYioIOIIqtk7vrXlJaDAOVyRtp81pf
Vi5zjFmckYyIQmrlYM2DWWGBYKbluyIFfSlzTyBdSZHvs84mgC1/R1RhdL/dP/8W
A1D9JBh5wbcoUhf215HrGkuOf1QyeWZFXVY2LMncBoFav3wFoYBKI1hSQJto9WL4
zLg38accyBXLHG4zWjMzkiC4NnKCx+g9GZGntMMPKe9M5Imfgm8RCV7aOCd72+pe
hw+leH8Pb8lXpKYOgK7XcTIVaF6Z9kMQB5pmtFKfbf8SMyE32mwVlbkgc/MxmnnL
Rky7yHkKwM9mvl8YZIg7MzJEdJ3k3gCN5Ky1H89RsmPvoYt/fPQlzvJ+04/htN9z
30huMkoKek/JQEMuzjrjeEOGzibdh4ritBrqQMsNkdxmLOZt2K/3r8r17uG4pHNP
NAMfhpX+aL2g5IZeViKrjOCOG2LhNmSybuIxvCUK4o+Ytxx5ViLM6Q1BgIVdKrvi
UfVC1jwrpmwKErXIQ3bJ+MVQHrM3obe3PTDtU12SQ4sVts9677z+q+3hJGnBg0cG
eNGleYPS/HbNMxdAilY9laZxYU/wbX9uVXZ2Sj7Rw2Pyx2B3MG4Wk+mfipZAagsp
frsrt1FVtw5dfftsaDgE1Mxt/OsEyM59eadQ634kzuMKNP34nD7p+m5n3R5vBVGg
oYi4E8jYB73H2LJtZJoQVn6I8nkl2eu5LPJOoyLYQsGqHUypb/FJl3o6BIoqQptx
9adBbPeP1pnIp8Iwx2fZufmPg17XPo5sSWUosEc8cmYtv1Sk7kHlAsUNjJwSS0X4
Vgy0NjHcR9ZkjRvb/f53StFLotxSKZeDEI/w3ZJcut5BmIXpPdLJFQPDos4BpiNp
N197mIcNHPUYKiXcEOsbMUxe7NwO53fkTZhupchvj6OvDFdp+kPzj1TXg4zUihwW
LbHqsNEQ9cvQc2lcSI5jljtBecv/fZuty3VLwnkW3vY0n95e9FbKUK3cBMX8AcQx
0hHSP464Q20Ms5pIiXPqXfZQ8sE+H7+Bmwe0psOULRz3uE4WGXhzI5LlfUvcxQIS
pf0ZNuSJalxCR2RS7aLwfBWVKo1ZvR5SVvLBZyoyI6gpuI4DBJeqwy6trvfjcoHB
EC8MC2U9jwtRJi2fU5Gzij8iiC+s/DbI6GwDli4Fl/0qQygpBGaVto0TAX8lMb/6
8TsoxK6e6/Ii1ZukuqUWIpFLgBiFeBrZZ9NhhVgNWWHCLNbi6Wj29cDQFjLzBU3T
d+hOnbJmUHs4DHTUcn2OCxlkOkczXJ+pL0Or66GCptUR/aM7THEwqSveCOhb9ekb
9GXoTTZSjchgx1TffTgC6hfQiEIE0zfbJE9ZFGsqCkADtGcGheUYnOA7lqvRQt3G
l7lSmIJTCTn4QW1uYirIRXipG0LjEgEnm6kFB6FeXI/6XaSBYA0nl+ZrrTxD/ebD
iR23/IjrqqxfkLgs9AC8Jg0H9aJt4sEUQExILI0g1TiB5STZ+rnGAFEniD9LlZNj
OodM73gJt4L7hZ04o/04ryahMxFgBVohycER7aVTTZ8EvclPV3M6M3cPeGxQg9Wt
1CpL6bT4U4cv4lOSvfTTJoHR64sme667WQ9aECDnI+UHzZLIdqvV9VdeBQQzayus
KJlGNtedWv+5+AJdiv0iLSwTSScR8hgNi2pi5hS5gjaDnSxNC351TCB5gmiLk9s3
kxPwRR77DD6jV2v9WJoL93QF051A5EMDEavcqytUAV+/fzzDXWO7ReKkZUAW0hxL
477yWIZ+Up+Gn5Z+Pkgx/rR4m3vYD3/+AUlegoh+R5Pxb/LjPboTRZpreVGOnvPv
IOmBM1TVwVD2zrmhQPG7ZFnrYy4UHPxFYhtbh62Nhf7luXAnIMmx+M+UKA5GwdxU
aHAcAgHV+MnG3i14uRe93Qg6G+QSoWlBQzqgVfG2K9E41qpzl3dJGtWDApaX9cBh
7hzVRecn1ijPVs1SMRR+HB08rnC6mFP96aMPE0SiHY9OyBvBftE2GP7HxrhiIui9
uvZzcY+C7cJSHLJ0OlSmdWhYTAnH0GNa/+SVGaxyerbij0An7Yge7EHoVFL4OmXR
f/QMBcsHrh/zFBJOBbJyXXKXSBODjmcBwoVc5blixcN/FfvZKEkc3jurUQgK7MoC
bK2PJYbYMQCAr9kPERZ0oO1JZ9SMDRkontkoVaVvTzTrOlDnbx8c7isjvi8WTBOD
kEg3cmdA5EZT7DRv6cixkJrc0vYIuP8QdkDq9ND3FCqYN6s1i3+O2jFrNd7n8DmO
W+M+wjzTAZ0Udfh4T2r1d9VJRQHUPKoJKOYk+Y12sP7v1hGkbKh9HY7r5+IMi219
m5SInpXc0CRDDXB63wwGEWqjrNzMJdafQmKopwGCJ6oefjcJZxiUDmOmw5jGlMjv
rYdaWpbFH58GX0I/knUg7j+NV142Q8xWEQlAWPjMKiyb6Fy7HeoV9LWt699LeFyR
ArlJeOd/j7kmUG8QWRnvhntxTlqxxMdtK0lHxI8JkkScKrdPXtudrp9A9HejXw4w
WDin4A9qTnXGa0OaVp7dFiWUj6767yQNknqboWq5iTWLiEDy+pyrmp61X78vC4b9
FoY3z+sbdyVvdKB5t3r+NrY/r+BuMMIuKleOBSvzcOVitukKQY2+N1veQtPWlggK
9i/5nzIbfT1XWyd4f7YDto48gWuUe8AySmMuSrcxj8jaewYqKYp0E4gw+zk92m45
KVbMAchzmEzBV3ReNZpQYpnsVsP+3OEONDbUZwLUNlDmuzPKIywvLZWjalpZaoQ1
S5kemy/vTEC+Vrz0MZPz+J4WxsT8EBlRj996qKQUL9yoINGTFAt/WCzMHBO0nu4Q
1MVFougbonBLd1f0VDNTHaAUuqgRwCXRILVgtaVKvNqN4TGeZ00AsFqDn9WxwVkQ
OQUfBP3rPiNP8wJFlg+LcH7IMqJamg8QqOTIHkrvNsY57u4WFZTmEHMSMTwwoDpw
fVb5U/Z9rbAMiCiooPbf2cVj6IyIUpH9RcDLmqoeLdf8ONMOGStGbwUq/U/OLf2/
loy5JZKI/FZ2ar4HNqrexxKthsyoHDTNenbXC05dAXpR1RZR4uHvQTCh05A3kUiS
4nNnlmlb3q/RWjzKWafllDR139bcIH0TkDcoTD9f0d5GKv8XV/CEhoV4XCSH9RXa
zsWjGPf7OJoIvTu1dZjWDOlrPnDXc3fGox2IpjUGb3gv5+QxjNBRwpxNv7xbN8Mn
tbWWWry3ExsizZZM9fLheZYWlMpOkUIpzBzuUHMn8O14MsXx8wpkFsiFPAEW+tV/
eOmvb0QZOwuXQtAWRGzjYgmPhTq9yc8x7jv3btNpQ+rKrbA5U/xFXvHsg+QPwQMO
i2jZXfy9fMOzg2Z6I5BToQHtK7fDYdKLFEmm5VT+tmNxqnLB085oaFFgmJU+aFlN
IykHtdslx31LWvBPnXMl0Ci2ipi/CHDrN9DIctnQ/MCTwjrIDC+lkMBBvBGW28RC
XV6T/F2WDbF9WyedyS+kHUQWx2GDQ0+7VE4zK9UoLA8ECozI0+SZ4e7zaZ85hX+N
mEJZDMOUcz/tkDdsBRt5Fr0q3MAi73QleaQzkjDdA+Ume++gUwbfhJ2VrSwCSAdl
7tw5t9tUvnlbEr8kUQA7ynB3ayzbABSyhB5KxLimJ/6QbvBSmuPdQbHMEh7IgzYH
RBo2lnh9a8fY7stptvsO6fhqjUQpRN73P5lpWWJm5Qgd5p9PtZEiF/NBW4FtIhx9
yOkW/xjzcJB+AILxq5aJ+MzlUxly8bkLFNV6/znrrmnLH3Nz5thKSBj1dBOt9TCB
SuPTeGppHIMXRl5K1PtJX2SBPPtZQYO/EzfaLQtDiyUof6nCNNxrVQLFrqiH/j+P
qZfBNxN7fc+uJyD76MqGpVtnNb8Cy/VlZhHkV9yZllfDXwb9IpGNBpsXldOKbaJY
hDuLL4CKKRx0aOTP3HLEgzTFsCGxTizCrQxxv8wWcEf+/9AZvIersOe0VnayoVja
KB51At49WaAnQortg30cLMleWlPaT7E+Vb5khSED5ZmQOmN/6GDxnwSwqEa1kyGN
ZPQKkIX2mtZAeleufuX7GxIfJOCXEExtbxSVAI1+3ZyS3fi/YdV9KxGWHQRrkjGg
X9iQbYDRBIw78gp5pNDvw5ncdxGOKMdXgYZA7zLyffT7brsYqlAf5pNnIeh7xmTI
K3RScFE4U/eH4nK1bYlNs1BSR0Mx7PIkq2+we3oLx2A3Ac5jw0+vwwGEdOBfBPTQ
nfb1n4JbvBZIV2M6ywLe3u5YDoQuUbn8gjn/Br2hHHvmLSG26wyyWzgQxQgEPDWP
wHyZebFXrb5aFOw3jdHfxRMG/237IAmfnIUlOYotJ9ZBGRhOfMZL2KbsRhXmzmb6
sprsVwHi+OA9k6RBzKQF1z0fnZYoAl2IYGAZc04QvVj8+YR3zNyp7bJEjZZYu+Vf
kymLWSPnXgJCfHswgX7wYzPiIvh+NO3dmK/Q4S8sJCHvdyw2kVktqmo9izFfJL3C
qOWuOgdbfSk/t7Ec4DU3AYYkpbzK6W7nemyJurOj2asX9+UdeSEf2yy6Lw7e4yah
Taq0zDSVHTPJMg+SYc0sZNTRYJZFXVvT8HwRTBjeoQxH4MQJLApKIUT4YsNzxd3A
rjmLaklX3RxMYNNwdmglUrEaE2Msj/1Ni8EfKdwu+EVRqXTAQY4kCFERvN6my0BM
saK8nKzL6j5DnhbmR0WTTUW36KsqfYL540RWkFf7ZAQ4FGP+C2oJ0l+V6wYTv4uB
I/hQaT3/csUH7j2HV/hF9p5fSLMiU3ex6smQdWdgsi6IVPMzMOGXCu6+g710+z5Y
6aRnLLe6nnzOu7Rq41AwDOrE9iAx3OmRHdGFeqRq20h4RuS+t98eR4p9o9OlP6VO
U5dm17IdtXGJm/Q93uttTMkzWjN6diGdHC2mZpBOpdQwNFpEywXQFOR5uZGcCBid
IcQNUao9lDbfSin2pFFY14AyOGkO5jgp+9/DiqBNaUPAehz9G3QovT96PlEjiZrf
MDFFYU66KW7qPWNzv9+AfRQM4yRBPLfnGMgajJKoKb90LXlBB4JxoF8P4mgzVtNG
zjndavxyF3ylnMM/SqBRp2VKfdami6A5dIPRzTQqgsbfPcwRrVxuIBmZaqv+bESe
B4cSuYkYszWDKAGVnrAM7RzbxrjzmvPZqu+uL4eLSKhV/jTZhlY3yHx8C1ezcFk+
hCvAfaOzIccmBXzfpYaQnPzWUjr9vrj+iEE1T5CgS+edRDV/yVxdSPOud5TTgBhC
Kb/HvKRydzBuDq6mngHZZEBQueBUoECldVJ1oKeS7mPaLTvpmVvU8rgPdGX/0ibK
A22wmtek9ShDC1mqRLsQeB8OVI7fI8GqvBoQnUzi1Fml3hCalXnrKh5+l8fGoC5s
V+JFIXw09DME+q2iXQzKN5TbLDQgrEFq9gPHJxuP7jer2UthUO40ap+eK9xQDVPl
gI2pm3xFGfTQgpVortP1ZD2XGUD9wZ+Zy3BjZb7Bm/y7q4pTw/a0NViWXz8D1xVz
XkYvQcge2IXZtyjzbpXUjMaKTeefql+MpbGBCM87tNimdJRr8puR9Lfb73ykFqUN
Uu1NLS4FXa5HynBcNQ1vcIOEowphZOkVAPGsLVIH4YKB2448NqwQOE4pl4EluUOD
9KcedsT8RSD0JQ5KpXt2SvvkIwFm7iebr2o76L1vUARp6sNeaIkzPrkZzp4foh7e
yhC4RcFkKVw5vUZD2AToyQItjLhVvJM84Dee6qfpcqOPWvz0ntpOeP/I5yhY8w+m
L73joxuHetNvhyW3ZVBQDkwAhOwCLire6Kk2VLJ9GSrun9aB0w5reBrIyLToKNk3
IBLcvteskpighabstD0UyuIOk27PiqcRKNtbX9TnHQYwMEUf5i9XWSBxhAedRh7v
puW6gMTJAEoPcFjvnonLE9MyhJPJllOQOsQWJ/Xkv+bCnvwWX/Wn18WLDQVA95uh
A2J04RNdydizb3QSndVjdNPeerTOz3zwthP+88g5GOEuT1u+qGH3hNgMo6fY4IbW
nycOmOudU4K16IHAYhTQIeXt3w4BN4z9QSaSnAS03whSmFYT3jNqpBL+QEWqHDCp
nCEQpo8loSURM3V4gM/3ziETTzmxLtmiba2ECkbz8sEQd0AJsgI2wekA2m10iQTl
zRzb/HNwOG6mS0riRwgIbNG70CCjK4P4LtB6NHMzlmcXkmX85mD2nK85NJNRDxav
ft8pPX9WkhdYvWJQRjToXMZ8EqT8uy2Bxz8QJgBGL110WLN0cTBOzNOLbA/hAXrU
96hMNPQunGgHtzhg6fSxXrRYoT7tYCtRrIdXf5IuBDK/5Yhe8zMGBS+yHq67coB6
h5CQGoM4ZZagdztblUAMyI3PEYRADuLwnf85KV+96XZWFYejFLtCk7CF/kej+/cH
3czG4O4SBlqtFgtmpPmEwhN6IQ722gn9ekZbDKH9rXXCsZWYSDIJUM5VA12fMMCC
wnmjQX10w5+SpODCRjeR7FLZMjm9qzzeNUPjDVjMvvbFtUfMDEr9NJEgXUjX+gYa
6LjHxOavH1lWy8dNDorE0yCzco8xQFdSto1vA/fkNhiMe2sxs0CigV1flq78WCTI
GpcyQ78NComras99F7YoserjiZVnu7TVY0EQZ+gkA7jGPjEae1Mq/NSEqnZLSnCm
qClBHBZxuudq8grrJ/+vITDBShp02f7nvx2ieMe8SBHOOk5aY3zoZXos9WWJ0Qp4
M7/MxLRgSYoC1BUyX9Z8KMAYQe/PPye6I4cnjYKtgGd6tki38tYb6dK1mKcnriiz
ZIUTHWc7JbaZuLnJZLK31LnMPARMw/3u4My4uHPR5gHl4wBq4BnEsgFRBjTCC8jp
n6GNHqIjz38f/uPRVK/emcO7PrC//+96jisQPJOTRTU5p0yW52dI0Z+umtVmKF8/
PGFo7KKHBEX2JrV6vWezZpgWX2g+KtVdWKwz/RJxGP9xsAQkTYgJeKIrBZ8eJRHm
SGGLx1gtCVKM6LfZjnDCPb3+imIVspuBLjjhu26k5TPmG39olGCq/nCevOQaq2Tc
yK47x/y3Wz8LnLn6d9AMThlPIfdoMZ+RieE6vZWMQltUCmUyZ8ypkc/EQCTOdOYl
/MWlseu+I2Sf9e5xiWmAhOXsJLOCLRcfc9gbZ8TvVUleT+PylApODfJ4tBj4Nirt
eiGp7dr3Q6sGDYjiI+HMFONPB1H4WZyte1pt5bno7QGu/DkWW/bwWglbRdWbvw5o
i+l40ZXlEJdEIswzp/IaLbW+87azdUyuoabAvsY8MhT53/uLM2JUasBFwTXoVTA5
9q2ecPsCfJMKjqhTbMpudI5m6LjA/bBy4Z1X5WwMUrmycbL+13nToOTYUOsdjlBv
WixsRCpHeyxFRoUwO40ng5kKB/JIg+3OTtt/0UR6c7RTw8vfQOZYWXjOLxM+flIa
UERTRukNZKPV3zz5lwOxqFoYz2k0qZY8kcuD4qk4onerRl1q7N/KFgzYMJb+NQkN
/p9sbrAfk6HuiIh9DvAJZ1Qsb/HHm1Pbqdw8NAFr3hqZ9fxo4GwFniqRbFAuK/us
fYg1ANBRcr9aQm5orGGFxsC0X2joLP/uIZ0LCpXA6twVZ06R/u/e/mEsGYunvQeN
uRDFHNgoBLLuLo0iA5YCql91V+5/0T9QalxNGab73xn5APYFVXhcTdECgbr40KNd
Hqwkv24MNPQFLSnZOqv6hif6T8v/10WYQwA309kuPJFxug4b4uSeeAP83AlF/bd4
mDIY1oenT54aXaDKr6JjjQOrtDbIZ9pwaS4DPRbX9RQs2BeBajG1x5nFP5CNf/0q
dtAWaZynifXmkRz0uAnwDIg8IxB9LsFcbFPk2denT1o9D1Rz23I5raaeASymzgY2
32BPV8OG4o7h9Zs0jeyJNvPExR/O1zA9HixDFBOnJSS/vMV3ZsDgVIKUZTBgFgZf
tZB1dS5LiNzrtRiRg6im8WMKdRWvl+9Osp/L2ETI0/DPhMgTKSsRQgN+kTEeMQ3/
Hylpitp/+4QByFfrDYWE5g8B7FrKhMLrK1iu0NByO9JswZOeGEw7+OPa/ZSxcfJF
Hb3RZTBggsHfBbPOhKlszS4NSrrOF9VevSCv/sc0ZbzOYO39WSchcCb3vsY85vCj
wj/EGc3in9cKQ7/2TmweBXh3FOe0xYy85MwgelsyIqceIgOfLY8IHD2vMMfzMp+2
YJ+i9/f+k4hYiwz7O4dyyxpidx5pI4S3TiRb7gvcb2puLRhH5D3ibclVbZfAVtUQ
zhN03DaE26bnKXCxRWOHOwnH3DOmSRzkFrzoBxqJ7fG8nja3/7jC00uLmX2FHDr/
dycyAauCKkTIpXdoA6z+9YVw8vQY/yXiSFXbEucbOmMUVdDGZVjJcBTk9QGKK8jV
iBXyvDz5Np2bOgRCF3A5EIcPgYwblTrSobGXqgdtHJT9F4CtNb3vIsUckzDEyWFB
js34yIfk9DGKHUNiFtp02Ntm597IV1u3r4gguBuvKNCV2E2u1dLxAvuICdz0cWRJ
ePJJbhx5/ZnEJWaFm8EwWgip14qosbMWgnpftQrcrSfq3ux+vK/mODtxTw4pxDHW
HUTVXWoCpSzyo6fFJfrtSbFISUUub3t8mdB7voYAXI9DdcYiK6mVRhXh5xFV+PyD
jY/vlSYQxV31eRxuMc0ZFneuD707UhfYxcJJBxTBNVudum3XsYFY+5/vqui3kPCY
np8W1u2p9Mm2OOMINgoisvcAxghpSMjXDuO4XUeIB3ZYFhHu83T82uROktcLh6UK
rjpDbMcJNzCWj7cAopT285JpeAk6YOOge1vdxWbx5EMSB49XLzRiraoMohi4GmP3
19RJHolkMazzlKWarbhrApanw/m+eDo6ZYZqL1yhwqbX2lY48cJWLoe20GUQlhto
4S4GjpuE1GlbupVLcTg5nxE5cCz3M431Fp/Vx0Alb7GI6WvJGV2bT5JF3ZR5TfZ9
XVgRXCrqE6iht96uPyMDxMOZMB1vp+AUDfr6ayk/0CzXSXetNWimElgAsihdKKm0
GA2SyAUaQfn1HAfu/h2UiB7OW8ROmC9L49J7x/Y0kCexLj2/C7Fqnwn7HWt5/W/F
3PLvLduxAVJptrMQ7d2mYY1g/QZE9o2RvtfC5vnNNV/ODA3JkqbB6EF8s3fPqJ+Z
sCVXiYUy7oMyuWs3mNwjU9spxrXgY9z9aeyHYgebRljG08FHOlTuAfLKOiXTP+Ca
lbNWvt7tyuPhJUS9K5mUl5595BuJQjfiaFuymhRH8GXXbbmGy1kyWgcDgO5KWp8y
wimDmf3adcjCcnopxyyuohu2wJb5Zb42WmeKYRRBLhjzBcIeZD5SdHMk0YJPb42K
AUip/Kz6KEyIgwAP6jSEjD8NIPjYdOweKrQc34YQQQ4STuglphbaomCoHXPAWg/1
QJA4pBxVz4YvWV2xYRRFSyk9LIiUEMdMD11ydBZqfCAz8j217yxGgz2QCGIvEp8q
w3SrmRb9iFr5ClVnMyJrrChg+v2iX3bNUUGf5oY+EaKGfb8T41Bmdp4dqPQMH7aH
NSBSLOE8p+fcvw1zoX5VYDqQx6e1w76TfUTEOUZltej52E4ngRlCtOfwatasMLWi
vXnryotRkTDGqLU3BUBzvKTuxYuQ73MaMMHeTic9mSvWTkRjVeSIJbSdbbfIN8LK
sXJQ1Y6//xlZetT4+EnoX+mS2gZg0cq3V7eJAdwV8DV5RRDIW1u0EQmh7Ot5AfHO
QHy1cmx5vkyMYS0oVWMYzhIjHW7uyOaSMPaR6LvULp8Fg64SMIe+x//X0aaxNfEF
BoF0lELCsKAktIlC1/55Zow6e8PmgF0jzTNcuCfb0AGiRFcaHl/i86rMLWgPQtpV
IUn5BqQULaCR7xAJpiGEc51cOMU2WgIdG4tSAKP57+Oqxc14Axzm9vUHVLpYVAIS
roVrm97Ud2uliOECg2RrQ+DKNVIL1l9PfZF1VX9rvBsvb6ONURUeFBC1kpGTAB/q
H03wylvTiH79+ItKe5GynaKjvWSWx+L7jew3Q/yM0XbNsL/jxD6ZEVPKp22FciII
SlY3htAeg/gAtpbexga3Li8kp6Ex5Z0QDzZqniO6YlIUS+05/jkoTrYjc06tey9E
pgc5kJM9pyJZ7mRLt5kwQW7CJk+6/S1MN9ra56oecbCBVqe8MwF/XQ4n99xhVMJ1
4j4yWw11BGOa21zbYnJasv0oaoWbV/uyH581P0H/QUYQFHdCALWBFrFn+hwtX3Ak
KKFcrDMZqRbvWe4mmBDypsUxjiIavp77yIPxSbWRxhJxozGuJdlW2LuYmgRzzVPT
gAZEDLFaNutj9/kYp34D9O5/tinyRFp4tOVP7sR0cQAcBZWyhMws2EUUqVC8pu0d
hYZr2aOjZG5uM9ecykmLXw/W9mlvebrpBZZ8n28w2v7NhlMv51qQGHXvaLgWoRKG
IO1q+BHlMAWFGferXNaT7sfImqnTuUnQy/QOGVeCg/y/0vScE0VGEzwPwqizv9VX
T1LmdRrB0EPiGEsW/YEZKC/Ow+t3UafynOs9ZrdbAQzh4aHURf0+BewG/SUagN6B
vXtAQpO+3yAx+y/b8mqjQ8wAeZRDhRhHZXMZVukTh4FnCDTi7w/wcFQtI4AS1oeU
SgPBky8O6WPpDQ82/jE1fmbWk1A2uOv+44umHunJb2eqwfq5+ywQ0vnDYTHwXfql
7qu9gaBW6OCz4GV0SeX6lIV6jGhvXHtM2r2BbLxGHMXdh/SwurA4sy4DbEOlLiT6
N8xJk+xfPPKmZAP5u3nhIEkXQtC1h8fjViPZRyxpc3QdFeZNIXroHnuMy8QXgLYh
ZJ0/Zn0LOIpAa+fynFqk3ZK9dninEFj/gYYUsyp+rljuLTajumsQKNJMP1EJZCWS
4j93+s5gbM/8iMm9ch5eM09lmLz5Jt3LMIWuRzvdk23jZ2LKN9NisNQSk3amxrs9
9rOpK78jLzqOEvHc+fh3d9vn95n+ixke/QqqdoPjQyCbk7xuGgOstxuAEQgDs3E8
h1pZpPr9BSV7iqMVdERIasNiXTwJCo29Or+2eFL67Em2iBdPagfUAckOmA9/1wKy
y5UVIIBJMiOK9edCD58BsXoUFEMjrfYPnw6qmd2WrGyheCi/oYrIvEaNWM6NkF7w
yJK8f1GVmvUjrkbE0L5ecIUONMsb0CsqIxALX8Zsz812wBgPnGrPpQbYUgtwiO0N
FXDey2bn7xrolHM3Uw5DLcXWPqY058m0NrnjPciO4C4aTUxdj3Wjl21X/ISfN3Wr
/X6WdRqbgDSn7WtG1pEUWnFTT+ZexZoBsigijOUe/I7vJSiFV7sdt4UTW8lbSASg
lbqpk5R3H3aqzO5E6b+4qamNsVeB7Om6/c5JvyUy0615C5NNa2UH8LbtGBnrbfSs
7B+O7Rl7G+PJP6IIfcC4WYB05LXnZb2QAFs/BAFhxC3qckL/vPEc5y4TGZNZb/1d
bKgJ9qBui5/iFNugAPwAHxQKM+Oiti+jNVYxuBUGuFoTEbq+xzrkJ3qelJb3z4bB
GFOhCsMfjvyEON2ZpZGdJguKXBll2yN+z99dD2wuIrHKmn1ktsC2EleJ5gwSbk32
iyqzSnMjUGJ5xfkE/+5sW8FaJX1vHHOGhoTyxGSZdOvJJ2ZAXsKnQC1JRReVp2Ui
5OEHSOT2WDVizv6aRtQNuNBivk6iz283Mbavqdy8eGPn/QOI4WzGDiygfYhcxnp0
agJI5zEz0a+dMIoDtLQOcT5kf0xicdheE4bBPRpfzAtBYze9RCAZj6ChhkzJtiEp
3DV7ya3S5qQWrmq8i91W4BkBWAj9gzTq7uqzG1AXXnRYCRwKi8ELCx8ndYx9zd91
HYOyQl5FuFIvQitSzr7uB5qQU1amncJKXFOfZMjACpjRcmfTOMR7h7zibJlGMcie
9kXBXHestCIGQu94a3Lm6b/eHxeJSG3WVr+RXSK+Z3K/w2qCTiFBLikL3sNDSXAh
ZKmor0X5M2E45goFlGR3v2+9X2z6y2siO8d4Pe6hP/HoDsbNO4kkdVTlZEYeGzrR
iGXJ1aN9HX2Q7fPBoINLnBgr22pjLGdMqXtYYKk7N/P9jWF4GYACyRBpIg+JhhFf
t58rXqUtzk49U+3Y3j61yUmE8IeNKNPxBktRPzrkK/dYFfBkrD11IW4+Uv2Lf5RM
p5X41MXfNPvxSs0S6UYRH0ruDOlLAqrs+NCX4CDlp7Si2gSqgU+T6HA6n0JAoICO
iXuK93LRFqceU1N47CoY0CpiMVuvVIln08puOCtudsSRLACsWIO7dmpYXHKKqAl7
9OvGXsbtjO/YRiNrUsqH9XeVFZ+Bz44iRsDDvWYTBnz5HrE2UgF76m9kw78dK68f
ku4oOwKR+/3XnJTn1q6P2ACadE9R7M/KuNR7rrF36dgustce6CvBQ9LcClDXDsau
R5+oDKRLr9u8/6CU2Vi9FS8xz8jOk7bXuGQUriS8E70L5Efl7IA0Qkz8em56MeCT
/fKjd4nSCXpfX3RgfurcEgMJU1VP6bokSpdA9oWOKGL4q/pOr5qS2G/fGrRPTY78
QAQohKsLcy9LJ1p49BcqY48FAd5LSSbzE2cM6YYqunrpRRqmtc46iW96ybfUEgmN
K3GskUuRgHoWHyjduZfptUGEHICBKIE52fbVUZWy303B4MivmzyfiZwOvkA8hsPg
26TVioget0eBe/WJqopRV2eWKmpr9dXpt5CzYY5vMMj23Ej+KUcGbyHHeBU0eRzD
G1mJ+OTUBAkYFpsVuniQTf1Useu+hJfAf1NVq5jPOU4n8Q0IErGJn467eIwDMzpQ
1BQOxK4/pXLxXbTxryusx0aXaH0h9ncYceWCugYlNaHG9n47RaTL+Agyf/fei19w
qLDXNEKn3cf5Hxb7sDjn1Tg96QJJh/+7bORn6uqk8R/nLsvZCNJDbBjWbzm4FIoc
OITwW9xnp3PHDgLXFQinovDL0koXQyVAQYU+vXCMjHiOf5waeHjFtJcTRXvparYM
6VUh1hg3YIrLvEn5nPJhB/X+2xVGGFTgNspgHOPM3jwzx6dLejKPv9/7xiWwi8eX
sFGixofcDMddXz5Nd6mtHb0/WffC0RIfWH6T56wIUwH8VwlV+xcM2tBRv1cj2CZW
VOadD4hqgbmRF1pvJxfL9TboRkcxWxaOHrakmt48JHJwagEXWuxP2YiXakpQzANP
ilj6CEI6SIlWvCjG1rdJaE1qaym7vlu6ISOyFd8pPO0MJKlxJC1ZfW9dNi8LfKS5
1GupA8qccGcAeSKZpwW7RkiMLp4KW3KJZY8jkCpgMdVVlsa7w39o1wScdc0aI9CN
Q/OUun3fmgSyxkSDX1VLL9CUSKtGOvIO8CI6RR0n86vq9L0csHbLDAYa2snBSIQB
YP9mxdn8Vt/wcbglnQxQ38PgvA33+qBptiJVoueXgpA323ZExClIIyFVysDYuTzV
/nyrvRR+pCH9EvA881H0JCaxQcu548QkW1KHUbxwfLItihtyJkv69PWBYvyHWoCg
rFzHYJ8asHsoE/TkdLRyQCDPDmSvgqdv1RTif5DaxUiQrFFvxA9AAkNJ+zzt962T
4M/eRx0ic3eMhGhL3mxjfu/J41xrHGZbiz0/BGHtrfY8W1UXf9x+bla3VFRgxr0T
rL5cN1p/nkTF4Vb6ekzPmcOCVuRT7GRmY3OBvy9TYtYvKgOYmwvSxW34l+HwDHBa
V6UprwtGaceFDwB7v8pHkQXUd1jgwpmrx2nGslaRup8m+Z4ThhHY7BSAVXHTGvtR
+K2encZis23QNMCq/QnzaFZ7x0fMexap12MohZDHcHcvXYWjKvXCYYUWj5FszCgE
ZTecxr+9gZ9/ViPurYpTdvPh5kUiG3qh87SZaicStFQfH9mQDhEYlHrQLeite9Wf
NHNz8UHvY1EI1MUuQFprt/Yma7TZaPwZMBxIJPCLre74OhRwINShffzG33+u8Qca
JD1tWVIhVVWAU2GBYOFWSxQKbx6Czg99BXd7t0s1XTclqR+5khrKiP4f4sqFYtaU
psg/f5sTE5ZadWIDSbAaFcT+LqcEAP6z/EUo1k3u88XJcLYLbw6tgEbiz5nw94FT
IRIuSQnp5sq0L6mX5BMBIiIQW2dqDQhZZRMrmzEuW8aYUBF7toiRlG7iBKbl1UY+
Vnu2GB9M4fS3i0UMtCd2Rn6VteZYY8FezUtTbOuOk5pw62y+ScDekC0KdJiwX/a0
adv1+VU0+dJl7TKwhoN922RqPH6iA70fS5dQ+A5p0HvxwIxOX/FWxIEKNMfw9x25
c7JG9QzZlk77Ii7FUIGb3yrlrMDEua2xmpa0pRy7QyvXRVS3gtp4sTIxrXyHXVz2
4ITaqLNYdMdN5zzVKed/LCldVpkDNDye0g82V+zIhYAcmMBibN4QFc/3zl1nz7PF
tWKF/eRBdTYTrpVgnhGCqnco89MVWNUrSqew9W3/utEMOYnbO15fRDEgCI8oDjDv
YmS+jXfOhFO0x3DLahXGwLgkAxt2HqnXYYrUWvlPB6Zcz8/p45HSrL35VDVreP9t
HnAkNc+rvpqbCRV2ke7OBp9X9trP0SK8Z7CVNaf4ZLW4tHxK82PAGw8WO330B+fb
XlRy3eb4OV33+IF3NWbyLRDrEfMmQOn7bGQaswcDU5swauLh6M0et6PEVk3dN9Gj
ZSRnWfdDKNErBQcHLUJSy9HEXlq7IbW1Oxm299mD2yGES3R7TS0BJMyHw1kedPSW
9YbsiGQT+l3RUT1s7A34wHn1yUGnxc+ra66q09NPhwyZxOLLOAclI09Gl9CA68nM
x/FqqcodT61atjlCiIZdUR8FsnK6xm2HunungFHT+MJ5jFGMx5V/1wWAZ1y/GNUZ
OqX6KOnpKmj8+WrAo694CuD3aicCUe1HyadW1B13N2aqegDGQwHmOXQyNaU4UDdK
XFz1e/+hSMigSl8LKkI6qaDjr5FCC3tl72yw7t9ZUlsh1hmMIF3A1tVSM4LJIFoe
L4nWCMJTkP2YhN/gqLlHjpxyi7ovoONjW6I9jbYVv5h/iCL2U7aI4bToN/lg4L+f
NGzl8QGcpObJauVCCTVdGs+X1ggkrP1jsQBrymyXlGbrFZMjzzoi5Y4Wj8sVDYiZ
kgeYRwgYC8L5vfA9Zthhcz2Mj5/x70QKdEm4hGXy3T9iwbwTYNdpoAJbB8yDFyZT
e6GDN4zw03eDAMt2Gl48tdpbTtKhE4/dZnq5GMp/ttfXRRmp1CCDCRt0s7SXmAGb
CbjXiPgHMLuruc7LzqITSdYIXxvXL7NHWX3k70BTJIEPDeOxjOy/fILYlpwEEz4a
BZaceye/af1MuI9Vo4R89XIe45BJ6AKBQX7pW4RyAbP8hVb84QTug9b5Zgp364Tj
gOQH/SVNdvNVVNUMffqDxydSkNP2GYX28kjK1SNdAqLip5/DUAU4eIEIgI8A/4Gm
od6J1oojGJvtAYDZ2o/1uWsV2SpDO7rycm9AtaDlXshtnfY0aos7swmuLBKjsvc2
LgufUWn9xz1D0mY+weB/eOVX/pWa99poLsFYCBvwaAh6sQuPSrMLK5QdmQeqhQoW
ZFdOGZecBcjolOAx8e+ZDViVtDBWOqrU6t4f40jU91deJATdHuqyy54mRiIDWgpj
OXBnBcLi07+/sHlvMDIq4HtOHnMn0iCa0MpbVn+7LiYhtQK/qGmFn/WAenUAC7RC
Jxo5Wu/sYLbP84kSIkIO/ncaplmJGFmQx7I2mkZts8TuZCGoj2gUjUh95pDZUqAx
/jZqQFEKxdchQKYiqw8tqPIMH7m/GwSgH+9mVY8LutgqjolOMlnq4nFxTD0lAQ5c
nDKy30x60Cy25cbeNMojzo+93j5PiFAZxRmk4N0Z6u+lG9KAKT5qYmlTcUywa5+3
UHck7SWjyBqXsZReRVe6YHArNFevn4rujzc95NEujxI5Q6nKtohNPzuuo6Rv7zHP
mcvjfleSHl/e/yjSVTy/t5KgAG4myyoNoceE1EVMsn+BbE5CN4xVEMKAIFhtjixz
KBvZezufWLR+59qCeGGA4Zd997ZYxkkDPrLbgiJOH/+3/mAjzve+SPia6upkqMit
lN1d9u9zRT2fp9qVmTqgQTrwFTKF0SMwNDq2f68yaOirBTwibEjsHbY1hdL/SXQU
ssHKs9PMFk+e+l+PbXcFMMQrNJfF3ZDycajnpJwujIGI0iqVUL6FPUISbEbDUcVG
PHCHryAdmN5zP/GkNG0vOfDtV0mR+Q5O+1iU681NuYpi8MhuuPOjOFY2IR4Jzayr
pmpN330xeqi54GO62sZE9/zMxNkml+rThAkIhGXP8+H+c/oF3wlWkcYezQoijUJJ
2AUoBIRLZCiKLd2Aotvr+IkDG7k1I/9j7q7ol2bLwIK0SwmNLb7Du+2GXPBr3eaB
i5plAp4SnELW11Te+LoCgxNMXRcf0RbOtXEu4OLuRMtVQfbsLt3E1L02zuFNfmYy
KOBPLD2AvCExEfpeMl+7QvW42bRLfLIa31TbOyZwzQC/Go46J3Wfo97VniJ2gq8j
KrjIGkkzTvzWXVDEY58M5o37GPPnJXziQ3l0Pt2Wx2dYtEk9bMYGsXyQ3mXBaNyt
ilwxeBaM3h7HF95rIPdPZF78Rvxx0jaV7xW7ZPq/eVRlTCy9V5RX3+qPRmqRzKgj
YN4+9YDwXV7PFokQ+mkSiadxNa+fTKoxEv7Wuszjtcf6mKIHAGNB4Jh1tyre74pX
Sp0bJA7lorILdU7AuPzx+oVmgR8yRT0CNqYaJFumejWeN3R7uf1VI6Gn/t3LnY9A
s9QXWAt4LO0/Uqmc6LzxS21lqegA/K/+b5XeeqMUg1+RL8xEu3cP41+DHzhfolID
r0oDat0z2IwKYGR7jLve5VvqMh0dlySSz4VTe84WNvVEO2uKQ9+ZqzBju2S7OUgr
KWTc9df4NZli4EYKKnUYbWHducD60pTuW4Y/jFqqsZPs9lqskYULysEdwIH3DhMq
AsTPAtQUuZvPvhNkWNeyZES3Y2C4PuTDfmKtBdsvQ9AmEZe/037fZzBZ+AedsoA7
BmWS8lU4gGcHqVLXAkY3jyJvkdI1bOrEZJYfsO2jurS0yavHwNGy3XCfOn7OT2eO
P6aEALJp2q+RSmle5zxtbKMAlBO77JOn2ceAzxeuEdWxl/hW9owIsBigS6/HpRsT
yWOH9MkVgfjNrQ8ZJLLUN6jWlhISTm/oTrIwx1OftMhSJdgGFwiGWafeSLJNEKDP
hl56t+xhjgaTMSBjCsTD29febyjc/pdMXGzlJXZ0WkS8vDuW9esDIuhyi4fe6IAH
ru8lG/TmK8tp0cnyTPRpdV7KgaXFDz/DvmkIskNFeL6/xKn2CQ0zY70+vMVpvgPP
XztkvtsEoWdkfFjweYxZigq04rxsSqAcYljrScKXNoLVHvnrjy2WLJBkand6TZaR
KpbjZNNjK84HuCSnghJouIi3aeShuN2hi0dFyN0V8Nk6Oxc0Ie2nAo5x8GyB3WAD
UmzFy/2pOtJQrTj1BP1teuiXLhdq4QbzwzId134sazC1ByQuUzwWgEQjhbpxW0zo
qdbQ4YFsMMvehabIEZS144yDWvWcaa1Zn0rT5r6dQjd/67jhIKqTSl9kDWHYwyld
wuwOnFpqPoEAQ6Vfs4RbSadyTPGs3paXj5phZuezUCJOfzeRC/rn0BaMDq7iwj92
GEripG2QvAjtCSZX2tCcdSPGZy4eJoXND3XgDquYDl7izje6VBgsiJE2FzIDSssX
YJyJSw/ziBXA1JUbd69DvTBMctgY8tKVR5MxajFfjCTAUS2uIIsx38XhZGRhL+FS
5WptE27YKbREBiE8uh2mSKnlqkjXoEL+lwKgV7jEurD5sPA91qOQD91egIs6sZDK
dAoyf9sa7TG6u1S1/1Yw1vX5WjTK5PNqPV1OwPWNS5x7O8ul3EUPXyBgJyKgM4R4
hum8h3eVsj818zDUgbwPE3JjNK5dcjvYcuEEfxaFCzsjs6+dgpHaaDrVbRQynTFy
oO8fc5tQTMKATlM0d4/87URuAqrpjyhwgH2mM9XKzzOwunC6B9uDGaxtqa/rQaHR
pYrK8fmr+NGtvXw6U+leu/pHKj7Sk7Y1EDQxqqiV1JttWJE68Hb27/b8CChkplZ5
HNXilXQXo6ThCVV7PmGy7N0YFRD5MnUBtACVgMrZCtz45JOsbJyE0NICS742Ebbt
rqGcrToQRbq5sA6kPHs5PLmvZrcJhGK3n3W+AdLVhcqC5uhBvHeOu2aJAqIGGBIT
4Zw8Zj+GKRDuGOEHMc9hpvCvvqI8vGdjqKSMKrT3LA5g2gaIVdB181rh5zBMT8A4
rjVzS88pGVTcw/wqBBw35dr6zRJ9+WprmyhI8iSKcHFhYBFpzKB06RLmjG4JM/ut
dIe77TppLNqIPlTrbVHr9JwRSdn5/KkZzWqivaKc4P4hK7caFi2I6kydHEP74a6m
4xfCNlLQHMQRfxX5E0aenNfg3R4Ri3S9N8YkuOz8/flgbKXOigl2XFYxRPkfTqAW
Vsf8ko79JxcC90Seu0871LAky3E9ZA6mCPubCF19YH046VE0H2EX8Vhdy2X43c+e
17GzvRsj5eF3C0w+B3D63zsKQXUcI22bH0Z0l8bvB8cOnrL7Y5DW/XSkTH/W218k
dJ/5kywbHqU874KuMym3tcTsSHRkncmSha+MzJXeewVIDQgXYXIasKFY+YpxRnRC
cyby76zmchQYRbOfyka8+9s5/zLJptK7wfb+nUGh3OfgjMGqkpl5Z1xCVKKQYZrS
K2UpTJj98gO4DIvw9d8HDOGc9iIf34Xv6EvJJm7cTvYpDh5xVSTywTu1yAK9x0bX
bRnwiT86cfJVporaeek6D07u7JcPPnwevLSV4XtnLaLAHJ9bTjdPwhO4ezK/Inpr
mF6KzQzyosDH74pMOTFc8Dlx6lkvTzebNxns/TW3klWpLFgiI6rw52JHKsIqk1g4
xrwjdJ/nx/ApnLitFR2LPlUmIDAgCOumdZQOYCJ2tJKAuw9OZL+CHnlag/eOKNgs
e7J1xFfOdd6R3SHebH8nY/rVdlE9FpfAeK08qrihCnKXxZWIb6wL76QX0EGihKnA
bpI1oLkNrLn233QKWnp0pe3lu3GfH2Q/qBjDFuk7yJiBZlxW9HY3slde1pPDxwWX
tj7OboGcVb66AB8eqsfrzozK/WCdg3oMEHFkC9H4AlLKnPJfBtK9588c8EnPDqlW
X7LWIDm4iiYPbSqCPP8gw1YZxuifJyZfJGZVhZtQ2pfBv9xkS1jVxO+yw4tWwy8O
rJUAfXrbeyHQk73GISkjLRRjnlEaZyYrOCplJXa0l7YVwfvcyqS88AnUidaXpibD
qsBRPkXPBG5xcjG+yLIAumZvjRB/dS8eeDlDC1jw/NwP/lwn5x1dG0yqGBqOisjG
c+mdOQUlvxFREuLlomDUtjr8G72BR6A4lciQ7lV3HMCNkUdeaEXXDBP2yTP2EYg6
qKkyFtRUoNqjSapCCYe4UDwROVl8oWULUQqlP2JvOHx/LxDZX1xSXWLMSUOk4A3M
x+t4uWgs1OE0Us52R2NiQI3vRUErAR1VymX0NUXREkqteMlSPsZDPFmEzKmxhCdF
`pragma protect end_protected

`endif // `ifndef _VSL_MM_SV_


