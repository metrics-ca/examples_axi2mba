//----------------------------------------------------------------------
/**
 * @file vf_xvip_data.sv
 * @brief Defines XVIP wrap log class.
 *
 * This file contains the following XVIP log related classes.
 * - XVIP wrap log class
 * - XVIP log class for scope
 */
/*
 * Copyright (C) 2009 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_XVIP_LOG_SV_
`define _VF_XVIP_LOG_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
T/mQXQcVSlz3Q83CAamzTaOCdVuG9t+exvJqjiJxzTrnw3OhKgijVgl2Fw9pQs4L
5pjAunwuad4x/vX5JhQ42VRa5EohzOqr4QKXXuOEn8maXfR3NzHSRR0xDaUUiWcc
oJ1tjKr66ldVJoLWctK51i2TPLErSA3RdEenaJaJvoSxqNy4P2AsHSeJD9ZJbHBo
ISTG5l7q007tzAjLqdyScsbPqs6/RTcljst5NrcRDzDZr4oOtn0Fu221IQUlCHqb
ybGgPNjzgTWOCa/kpQ27uJrwXDegfe6yUcl9JgE7whaaprx8tsldUHox4YSmX/mZ
TfzeOTFmZ7r81x0NoPnfMw==
`pragma protect data_block
4GjVs8wyz/GxxPWSI6RwvvRu8rECx3iZmrmEgUwcibz+el9kTJnZkCIfJsru6o3E
/ctAqOjshIc9mT9irojivm4hzf3xzEaEDpSxXkz93nBytQ3RGv3bjhvGgL/mcaiR
HU+26hTgKlbuJNq2sFb1bKfX0IqWHC6elA+jd9PAZWyL32CvSqTo1p7Uf36vR0N8
QKV85G8l1KfvaGiPG4UV5JMJiiOcZIj5MxBNAETEoj84wQ43R1scnuTYhQFd2vu0
Swge1uxZmhPJ4CESBvRxxrrNUrRThAKlPthXUUEGlW6mkVIBCsLljvrmA7/YkZzX
SKDA4nVE/uIlhdvnOnQ23ZX7Hq/DUgqWH0NNra3XlGq9N0EvNcMdIPtOt6Pos+j4
ahMc6NnjAetR4N1YXeloYIOffX7iggXRC+lE6pj5Ww7WjxIzZKC++aiSWHR7JHZM
OYrdxQWH1+eru0uSruFdRjeUqWk26nQk0L7ZUjeloXKbZLqydMW7m9IMck9nOHh5
5I5SxWeLS3Qtkr2tTPkpVGDoR4BQ0sJHej9gdmzXTnaORCFXHFlJbz2+BYshrVt7
gzSQmZRIcHd33eISARRB38wr8vG8/Rm0aDpwIYjxRm+bhtch7vMYG5PxDFIoMRxU
feteuGxWdk+kvSMdUeyxnodX7ExWhQCNxEbMQAlrsUPQi+VtLrwvIssjBAXWdqBs
iJoiuLj3rGGQNQf6RnzvLB9snuxDwxuTc/xZ7KRLOJuj7gFzVMrMiX8tpkCfxHAA
XROiOsXwtKD17OjP4fvhsugAlS7eb+D3N4t1xdivDCA/I/+QreVvtrmCieAStBVL
9ChWaY4Vi0I+wUyWblL+gPDwcGVqnAJrPyMqgmnaQMOXle/UrckQTn5Ric/NkA7f
81DX/87ADzmfJ6IgXOrGaUMcVhiNMilw9DNiefaef063UwthaKlChgPfY4KBpnF/
CyzO/ytXNNrAhZycHPul67eucYo+NEjI82VaHceTJqPro+k/ZKfFx8ZnGPU9NLdE
rjbrRWdJaLQqzZTcSdMLhisi8eV5YSyoZp2Ctjceczk1QLGRavglRGstrElFPOdw
heOKN6MfswkJ3S6XRiTyQRrtxCR86PgfKCLfu+B3zE+pcaCAREmqmisESMa4SQWD
jmDa9++UixKB+1aKIqs1/9NHouoznCRpxLIY9ase9RzjtGL0jeLiSEyWaBaki3X4
5/QWqVQMXEVfLkCpMShO9ZDI7WmANGtY/o02FqqEB2yZWYYXMRyZEKvpmgvcT7KL
7sjuxo3eeSetLrCRyTLCYx0kbu3d2o7w801Ae8UnJOkC7wLofpAuygpEeJaoL3Pz
TJnRWIJWQv78iySYT8yJQGOsaSbmnRglovJwOi9H7KMb+DsJoYxnLSfTHwhdemLC
6vmkl5gNYagxLTUDFlx1JjzsQjIBGvmef2dwJmQ4fQMIuA/yZQKZYh6uvKHMBJFF
Vq3kOvRRCZylz6DMLhLAGvtBTm4bV9XUOf3D1lH5pld1AWPmCHmiC20kEn3VSBkf
IfflnpcV7T9227sEz01HchurRfSyeIqeoLsbGKFqJsm7xvtmABq31r8K6GYtiZDp
FArEQPWl0VeVKTkdAZPxTqEh6k/tH6iteODgR2y4uVMnAd08ks0ThJT3urfMWUxF
6dZB2O8zdU60R/Pi++GnRHh/bsjvdmPORp71e3mavfkaqgK/4tmGzSI3piLLwDmb
Monb+P0l190YYAcYqy/WIDg5zHJn19KaaSZH9ImZxCXrddjharWYOlCOAW8Ex9dR
C8YmgPoNILd9IwQGvhFXjcC85l8jruxD8tloaLIwebBX7za+u0Et/P490v7P7foK
2jbBzX7ZrFnCEaMPzZPNBIQmQB8hndvnKQJyzUg10UsmxVtbIv8oAG8qnK4ziNrA
rgBw6WCnDDsEErt6+yh5ja+izjk6kYi8g9jwuieJKE24sGpNd6C9adWwDoi6mJWN
9GVqEaoK+2jbC2FUya1B8aV1TePIJS6+mHrkyJjw2+SCLRROfGzshkoA1+j97Crc
5ZFn08XrNUS2o9gnoCtq6fXQN9AtOh7V8wI/XrEUFK2cFkxPP7sQdLyk+LV8D/pn
E9Z4UDj6T7q17OXrkc+2XGGpXdwcVDMON5ncJK8NcPR1ocvtbKJAj2yMsu5/w9Wy
bNVq8HRFR28Am/0h4zNRTaO2fvVQ46KY9ldAFeazL0YD79gkUeRlpVgdh6ucpEBH
G97RETisBD7Cz6I/aAUbxfEVvhsJt3y5bjO1MtkUIuNVerXDcJWlJO8pcT6ntZj3
jtRmdfrA1KSsjx7G19WG5Y03Npt+DN0vp4rLXg5wTdpaPMW/4FoGrvsiaWKhKpaM
jW/ss/iDTR6LJb5Y/fT/3HgwO8x8oFQdrEpW3rqJ8sxf6kpJ5u6e/YGtkYEEb60C
K2e6qWxg4Q5j3upHh1/Q6vfiS4HKuOMqxNMX0SaakzHhVnac/953CkqYrGbUjqDm
/sHQ6dNmgvYAZmWrv1htNWkAlz59famqNHeC27nqt+YygSSVlXtDMtiGXLCHKr+x
f4wH6WnDoJQ+Glfkp0pcTQJQUf/xXv3T/w1XaACg6n9TsuaQaqFYVzEAbhYt1KG5
aXCVgAuRQ8p1t2ObcqyV0gtUrvFYxWzQrdbtamaJD7RmeyDwBPz4ga1TNzmrV//f
L+nXcM2LpRh9mRB4FFStZQqwZXWgtZskdUBG2rV8AybMAJkin9dwCMAz9jbXYD3u
r0Nezzf8Ga2A5SmQIdJ1QuZIEdkYC4oAp96QEeLXMpCDk5nTiyqU2IYi+5rJNTE4
sCcGikm2MIwE1e7YtyEYczkp9m324Gr4fGeEs1qYvrPC/q6clVVfYKsWm4pVGAMq
tEkzoicfybaRXQt/Op6+YVmuc8LsVcXiYlU7mSfLXss9FN3qY5HkE1IDD3A2g9kr
ivNOWHqB5X7RqDJGolKNHSfimOx2MJYWw9GiF56IabGaeGVH/NSO192u2V2F0ACP
F3+FWz+jD+w28D2kT46cCl1Uo/piwf20jweoHY1QNJtbh5eeDpMVg52PXVUp5cWr
wZ96wNVMlTFSslTBXWs6mB9JqryrkuogZWpVs6+r+5DcwxjdCTH3FOx/cOHOhaTc
3wHWo9/75/kGFivwfd/2PUkeCE4s8QFTHTq8QW/FwRJmPSf77W1ddt4oAu6GAZGw
yAeZVeDO4GfznDSZE++tDyF5AxG0hGNkD2fMLws9IBKd7SDRMXiLFc2Crxi+S8WI
syV+aD3ydcx32pNtLH6jq22aHQ3EO/heQJigF/AaSMgfQnjueZ5isv8NreQpgmsQ
eEX+Yqzr/098DyexxgvHFT3XUdCBwmTmTx63refqm7kKeLHpyXiIKO9eBBpK9QqA
i7SGdK5PPFE64FhxxQD/SvRKHhPyyTE3xc8hEaXICLzBhQETqZxIXW0aRC83my5o
V6wG427/5uyw5lv+RMDNJVxn3Q6h9W1vrUOfURwP+52p/ig47LMUrU5SZWymBS+8
7vvOWSMpGeflt/Kntua/xLWfFyhrXSKBd7DWba1ZjPryAGPjSkhMa3TiJT5D9SL8
UMVq2zZXp1ZKBc+Ihfte/0HM0W0tAa3VeExL4i2H8E41R3EPLxPBO5XIReeuhKeh
3uvFOdwssXUVFiW2W/K5Qyu2+Q3V4NNybScnJGCkqCmZeVsKAZ7o+/mdyOF8BSZu
Ba+u++psvRXtXjJzzipPcgZJrdKmExdS7qbvk/+lYOnPN4k+wtKi+zcPkR+r5/QV
lNAUhqQczu5ShmxU4CCN1uVumdw1/6aWZ3mISlDNX+b9UZE8n5ujWjjZvDQzs1cB
rZymteTd5RkHpmekJ4CG+b5Sg4GBs5Q9bA1Qn8lBbbo8Ajia27XroIMYgs4GylTL
6TMjEpGrl35Jc6J4nkOODpUl0oKIRkR6PDwT8WHnztY5XZQOnvOBD2punEOudWqA
E/nAFf+Wf6zdigqblytW8M/X63MkJqXdDXUvAOIPHmh46s6R7yp/9ogdWWVOm6+t
klDgUwkBbkHg7mo4jd0342Eh5HTm3Q5f87UIESPOu60qb0t1WX/b0YaVbA0Q2nJO
p71DRTkbH1sffb+7XoDjZBkjSMb3RBO0L+r609qmyHSn+IkLOzpknlDUfpZ6uoz+
w4FTt7Kgno0a/dnEIi40sY6aDgxhApzCNqJ1b5sWuEB57GIyNAPJnsuG6MmaNxF/
RrnntpWnbs/FqvCUPHDfXS1f1jxReKFiEt7sonFkA4qpf/IzAZE7NI+JIOFW9lRh
pWfnx3A7NrSnixtkfxZ4MvBJTYkhpLFPp8Hhd+incD668f1DAi1PAqEeGDE4xuHX
PkDW0uMag/YjGMJdAAD6DKtNMcLOI8OfvqiJNaAJx1DxIk9qFe9KMPSuLAxQI2HE
quq1pT0R3SnMdfZFUvTmVavj8hkZaBjmQyCPlAcw12gqLV0nf+LXBSSi0PO5mkfz
Ixdk5+qOoECHksSDw9mwCB/tqW6r1QhXqsmw1CU1BimkoDAiiR/IcctDnOULcd+q
al/VV93IJdwxRCzZ38/DJRYH9i7SvFWvmGu8ggAujSivjyehlRuzNs0YptaNo71c
HddUHx03XukBT4QAL2azU0iNbTIKD1JB5I5aT+X35dK6TUlaN3vsra46ZOWQwIaz
a5H/MO8UQ669SC8Wi7dj1lWsvVQehtNbwTXtdQdC1PLfy9WmHgojRSgNUAtr6JZb
oR200gQC/rt60O8r744EpQA8KBHHs7ZX99ftzF6++mhtkSmGYB4a/JCzYMZmMDEj
mmcCziCVvD6p8gs0GTAnhRJTH7VUGy9dl92XIxa2edx6ZZ1LfnBUGiTfZEzh805o
wktDEwumqZvVl1LE+rgUNDAWpVIQ3Q8STrDaJv/uHl3Bx89PhDui+PIcCq2a5b1M
suaH0NlRDSxNaM8FmJwB3LtBFjgHk5NfQmIAkjkYdvGfE2fuKbIyssZBkejEZ7mh
vEvhZ0p6aqOuX8TwEhZvQzBLuNvz/y6fKbJ8TiToNJiTp6lTOQEYcHSY8XX6lKsl
N+rhDwMwhtJvAyERsRi2Q5yMzZ/2C+o07UNmKN4qixhkfacmgA7E3yCjTkzHt/gH
/aeRd3ayf+RB5NSJhYVRxUpIKr9op3IoR8dRPLb+R7+0QfcOgG6KnBGEuhB2S7Ml
fSJymtBR0+cDBCN6iV662plIxAb8D+ERlXsofzZFD8bSN7095vaDBM3qEHbXqRE3
6hvHkI3ZLuVqAmTqCZP79K/x8of4HJY9HjeGjIetQfU5cTwTm06tLP6uRgvXsMFZ
37GCw7NSEjP/WSH2JULs9Zs4mHXAA4zc4erQ48pu6JuqDMX7Sb+vI2n5d7fhELOE
T7Kjlyrpu1b/PLzJs9U0oR+YX8wX0NVxLCazv1GBH+zz39iXoN75eJ3LX6HU7u/L
j+lfxYCOXj79fI7BOJOhi5edFzxjoJFxDdkstgwFksMZd4Bcym9bkwErvpQv8I8C
L67HZ1fHAKjvfeQBkWs1PYBSLXRsfQf+3V1wlPIP6B+fsP93I+ss/BpaaaEGoC4x
R8a6LgBeC4G66GOCXKs08jNfWvtQAh8p2NDiU7m2+6A3nT2XtnhrYKO7LJyZiTOG
rGdMpDo1/wqBASA/YuLrakC/2PV3o/tTObwVazA8sQe8T7TV5Crw8C/SzxdExidP
JIUHdSNtSg/PMAAd2S5NI2F03yqWlMslJqRtpz5aA8u1C8o+aWZ/iKynxXEHbVqL
hgZcmy1GhZ+auumlhjZGemwKEvQGwg6aL2om8Ym3K5RoIrMORKsUJ6C3TO9oeb1t
wfJsnrFLIa5FoKwypG5VyBqsbQBczi73Um5CzR4gNAZ9Vl8u41q7CTp1natM5pnh
Tv43unJyK0yU755jIDvIxcLzeGHHJ+gaDhmInlZOUMxjKU7QIlhQ1NporBsbA8Ci
CXTXoOkNMP3ziZVRRS6sVN8G2sNHY8NtFdQvD2IIQEIcmj9TVif7rSO6lslTAnlc
oMZ0MdDpxLlUzWefd/+8Iy20Eu6k03f3CHl328/4icnOyJHT/sfclDteOfVFMMnL
hphjhQQK4Fa3J4UAcwNRuSmfA/X9kBC2ICvhQbc1C2Sj2i2OY51Vv6rQRgxAuTu1
qAJnW2YaX2d8e9P72/OJclegJWsEXmG2zi0T6bJkA/KOQvd6wo2mqq4jIhQQ8/tS
CWojgsruHB2gjHwc3L7KNUnPZVzSn2rnLTn5zstW1gfKkhUpCjSoU8gCiiK6XJWv
61LxLd09U+iO6U3WyeWiuTPVnNMcZclrnMNNSNmxgfvDQplyF2g7oVnoNn27eAh8
9rd/A7/B9RbSLdVjLojpdMH40gisGNFL5urEYVntPryjnPilwAERyASqUyfVPa+S
+tC1fWk0YaRVcTaRJLDb0XMMrw8ApHchEt1DxAkbGCNwPILKFrBuWiD7TSMkJAty
+sWinprm6dU3lVFO9dAJcCJgF7iQBIwGo5JqvgDWwdQXytxwtZTvcrUkIoquMn4S
6z8Dn4kFkz8XDVM3iqIVr1wGfZGQZi/YJHf/nSXdzn3jUhQ10AN3lU8zdtghYCuC
xDFv6bokEXOlIXmVRhY/mL3XdKQMIetiqrCWKLRLOCNiFADDOHjQrhAPOcPNmHeV
Emeje1GTK4S3t2hiaSQc4/O3qJxciTl0pVXy4PSWJX26oyhSyE+g51/iwJziHxny
roKEc2dGHaYvc0sGIXiU0iu1gcSreqlatb5FKlBdye9rlNLVLcDlF8+FPG1STM6d
Fms7ySCV/hqxrGKQeLuoyPFZyMv/pC0mRChhMahpwq/q2gAJJfZOhHlPDCT6kVNE
FjybOf4vjw99js+EuHsx+DrM6cKq9ngrK2P8i0hZ1ZiOu/QfAZ8ClK2W2PO/37Op
SAKsv0APWo/kYMQAx4BG6F4Jo9IxUYreyWXvvwSmNoo8i6x/iShyKTrmO+q6cRcU
8IbuN9hMpq/oXu3PuZ0+Rgcns3otiwEnxPm6sci6XGr9Ce5i8iZUUJ/v6VqURoy/
0cC5Mev821s2wLxLN2c/hN8amPWnefWd3yjm0vP54f29XVsaCrwu1JDRpUd95OSd
ks9uA75x8btLI2U8FwVtEMNEDoUbsW127gEc14SNdAP6OnA6cU1anTtvRQJX+0jR
51UD+RO7NHk8WJjDM9UkGdt+tXS+d0BLUQzDJ8lt9ApTlK+bJmOtw/Ge7RClPUc/
FjHsnxxy4N5Aqb+Ud3xdtsIcr5ayiG5R5nEDr4O2JjyNOZ0p8Io71RqRcPcatus/
p7uZ729Bc3Tfx4h+AT+DdD8AmZy5NG6Zc4/x2mVOlW2G7wWZ+ARHJj5KkJWOR5MU
0e+BBHwTafbrLqANkl0T4jXsgxwRBpimShBGJkCDXn4aerVb2FO/YJKAt1fOYbt3
7H/Ftw+7cLXI6pN2YFAd/CFz8dka0/He9fm2iynoR4k98AzI/9Bf5kvlk9cbS336
VulNHskGumCzLTFNuE0UU67V8qeMddMrUoXVHnfo6onxcwCsTIy7LSZFlf1eQo7h
vTahf3uFVROefGixLvLijrk8EZXou2s4oO656FmuSPWJyq+CUHzWj21GeDF+Bwax
L4La3AF9Q+mcbhedo8LRoPibaDussjg1+T2BeON/GmhrpsrQbl3M0tyfOcFc4MzR
Y2Z2gjSVunyDAegRy6yOy+Jca2uGx3KWwCXIFitrEHOgrd5vp4dv5H9KKirihuKu
OOQXbxh0itQR3If8fk0VoWbESJrtnJcpetzxwuOxapEFL3vnZ9bxma08novz9NM+
EGlmVY/tNgZ//ma5WBQvHoQ7RmIXHRpjcRCsxqm69DgwOrZXgXIJ1uWAKbb9PTQk
Q4LNZoz51Xa9EUlHXOO1D/5SNS7r82IPg8ObO1P+4EJnqy45D+1bCZKo/MBneBac
rEmwxmfYANQ3X/Ew9r6sm58oT8MCQazvnafeeZl5dkHN2wVSUwNDPDLvxdKSQ8f1
FTZha9+9mMlXKeC26r02ADF+tLV3tOV90VkVLYrUCAIueVWC1cwyFg6KFHCrKwOC
cc5s8xmWh7FV2CbM3WzURcurQOMh5PsE6wytLFuGKfKy2apCd+yv9Uq6H0hfjMYl
BeOUOoTy4KaHlEsdG80LLzI5fqOEnhgU78mfmBXQJdnU7ppCDrkxVKaawf/z99XH
+Dy8Sd7xIQ5bSVH4h5g/afszwrQxEUOCvPtV4AhCg90P/OShUSyq4wkC6dZY6Ymi
b6U/jNdbUc86k6VU9l4Useqp3XvMpve5uHnfjG3+ZcCX3aPlWFh+/D/zCiKAV644
gulSQ9RxHq1LOOpJOZbRX+tm/0FNyFPz7GvQetL7xI0CCqlryWFm+hwDYw17c/Kp
IcwcLnDX9LBIsjht5sBOAgjGI8MO0dcVk9/anmP6rHAq4OsY4ttdwmtMlNY25n4o
lnWRp56RhK6bDqUBk3NWBjvKbLTbh/n4ZTfv9DX+oYj++4yZriyG9e5G3ArSPTnQ
8gDWO4vQPWBO6CmW5rBfopl0YR7wTf5AsqOMCvBqfreb/ug4wwqBb/uju3PcCuLN
g5HTnw9IDoR2zlQMheiufmgbUwLHLqJ5qaY62jXwxntqI0H7rnpS2JXCyD0ypJgX
/1r6qlAEzNfiM6lTSHQIPjIfZA0Ye5euZOzyRXzey7a936DennRqqRqqjurocidK
x7VP5Fvhuskwu1L6oVbXhwMETvGo/kjkIFxnLTsN24wJVeiAXAr21DEQ6wOpANBf
`pragma protect end_protected

`endif // `ifndef _VF_XVIP_LOG_SV_


