//----------------------------------------------------------------------
/**
 * @file vsl_sbe.sv
 * @brief Defines VSL scoreboard entry class.
 *
 * This file contains the following VSL scoreboard entry related classes.
 * - VSL scoreboard entry class
 * - VSL scoreboard entry queue class
 * - VSL scoreboard entry queue array class
 */
/*
 * Copyright (C) 2007-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_SBE_SV_
`define _VSL_SBE_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
nLfigR7Z7pq9uNQtX4dR61nSPAbKBMGftTy6RAPSlK0GmIeJ1BNjc1Nc7YaiYSD7
+/uf2/fps4e+h5PMZH4zfw9QRoybdD63Gl7Njv/rAg/xtDBBR3T+cbCLj1Obejr9
2RN/zfnhiM43xKGGPr6bZeEBgHwxqeWGmRjdC28Y+KDPsYLevpPmH1dY8Jio53Dc
ggiFGcB0C+KNx0bcAQVI7iSxFN3rquIi94q0BOLe1JplRGCUi+PrvrlmkU81WX13
AUdPlvC/s/vQpgJ8xF7zcz/2tvPiInqd5hgu9t3DLVF2C/tWVT3GB4TyC4YZKVXQ
VmiayKRikL0viYaQWLeLAA==
`pragma protect data_block
rc+eBqHcxkPQJTrYr2JRfSBpISJXZfCgo+gneJPkphmXdybNvQqjUf5St7k7yBvi
BDxLrFLDMOLw/XJcXTlhzeD3jzr8B8cwuKB7RVVGOrKnRPR7L0PsJZKigTJuWcHz
WJ9REK5BcTkXMyqksQEbKOnmhYOvQ9iaPu/TW3k1M4u9zlcXR0lRaSffcdVlKRRn
6q0tLibZq3RLFUOvtShZ6IN9u/2li/rrrBeJ0BjZXe7k5EjvinDrJjLkIrr8WRuG
l84ZdOx4hJN+N+TsIOjfl93t5q2kZkmJcvdEQzlEQ0bRyVyF4rV69fYfEgOz0g6S
Tw9TWK4QD1Xsic5ZdoCyuklB87l3D3k+qnehFPo4iR5+6x7AjSFckfoi8k3cu2KT
4BCdwimGNvgiFoEYlFhNAa7HvnmOVeW65NhZxtJOm+/EmJJYTi36siHHvRddl3EV
sEdRHY8hefX5nkBTh3jxRsC88cl81Ybhv/fScAg85ETEaCcguvZAzVxdmr5MN0Ty
CRk2urJBm89E0DQzdwXi0CDCAxEbzSUmt0UU03p4RJxg5QYEBP+wZ8Jr//w5vke6
X0agWQ2YcrXP2wb5dAwUpWq6W/fsyvLP1bdtJCVPyDkoaeyw7o93kNWSKfMdOSGv
OqDasD2w7afo7t8qTeVXkMdNLgu2yew/yqdX0+OV/ir3/BR2EW6C7hm4tFZWgMpW
sNqy0uX14e5au+NDq4rQ7BVF+sk4NB8EPKicJaWRsO8sz1I1F4kq3+00+pSwm5+N
cO5JRGuj2jEKHBXzXQgDkcWETiT00hk6uSum3ZXdbrT2vhtwBv2qdTILfu8qjguN
idPGcnqXeaJg7tNUSBHk3CTr7fS3s1Adn66oVI+vujLOAJwWAtY8lEI7FxYUnQrD
BXnPpS5bDtOoXhe2Sxr3Vp5Zrzgcjs6kmC2Er/2NGGvDDsIv0PknJJ/+kgPE5H0O
ZB7v/1mTvD8Iln14oKtr7cU5T4/at4YSxDMvjuBEkn3yjwcS+P2d1LjktdO15klG
1TE5Ps1dzKTdkzDdRGOymoME9pEfuy7pL+v8ZqJPBc7rbIJ1FlLMxecOf4cXALvE
AWU5hoUDANe32dy+bJINw9nDMZMl8LhGG1iJYfP0bjJupc9WkNRNctYzy7JabQs3
ZavakGFNT/RcSAg6LUBU8lhYuwefxHAbA3bA/iu5zKZEzRLh29Omb0t3VA8z5X2b
aYEsIfg/LhqWp0xc8BNmxYTDZqyCcHwUjfvoYdHelpf91EX6zepoExuFiLHa/c54
MhNqXrJ8KnZ4VKSPoYNA8yepcSloeDlxcKYQC9CU+I9AOJLI1AOg1uPmAu1egeIZ
SZ4NGkA6AKvQPmvPVfD49bWdBJL8YLzrWY4GdM8M8gdJuHF0LlGsYSPmEhjf4AwJ
t3lLljxQTlhUmFwFLtHD0y0Fe0qZc5DqxxiWlFt2It31rxgwTGcg8/mP5VlPON2a
6m4NpYz48indXuDXtwstt4KuPpJ+7OQEzhKPbvJZHJX5ckfbcRQEishfoead2Ccj
dlHQ0S8Jxi59d9djQAm+aHNspI2HD+GtINyaM3ltGNYhFCprzpFsOA7u0rSS1bOz
iKXRskB6AA1GdpbqcIkKLmK//ifjB0oKUjtTa26WjK+EAcgSDaJq3AFYxQdGZQo0
mj+muXwM3zacVUD+FIyIR3HqGJL67gbcdjL/SwXGQosGwci1TOOR6HoR7/Xlfb//
bKRek6WZ3PydN1RyoRWw0YyGMSLhoov8r4Ql/8npezFF0LO89xIh0oEhZncsog9p
SvDQD+XRXPqLvFHAf+BUw5QI9Kyyob9dYHs3oC1QfF1srWtE5iXBh4miKgaBpM+v
yz4j8L3pDMFSqQnbJCGr9NkSAWsbkXgTCQzmiDPEV7KBN7a8Dfc+4KByU9k39O+f
uVArUJpbk71gcYRi27ZzSTZfbwzDBMXRg5CrsQi8gP7uMJDHrLcTKNqVMDBsrj8G
K570z+xdv1VdTDUbKbs/Vd6pmAm/7owaEDEO96Ui8JZj+bI+w3QeVbhgTjRBrCHJ
NNlA3DN44ooUhaVRgjIq3n9i8Cl7lQAVHTzw1IbFNHMxkQf2RMRc/r6+2UaRvIch
h8scDd0sQRMWOtlfU7rT1eURXTDbh1dtJNSWDzDpcfY2yVXbOD275Z33XKN0k9Dj
HAQrANUSRblAFNTlSD1If6flYjup0MvdiyyIlbhPnDjWXn0ZXakr8geF9IhR1tIw
n2qU35RxMmaF5dOM2FBguBAOkAo77v62LJIB5FBo3s/zKngBCxNFdGKfskYswnQb
radQCs7FgWL+yIJlouQSWIQUrrWAdamdkiJBvRbpNUGGjav9xFwhYrPjf6Z6wbT6
k0r96WQ2EDWYaLj39Lsf4v0gj6ptA4GoCktmPeFOXOQYQhyyJclsI3rgluu5RbD/
mIruwpkpc/Hmjpram8CVb9PTqEXM9PKdNbqVRrb6+s3uWCq+JHcTE26HFjpt/OwX
rABhClf1F68lmlOMHmx8muiyR9xcfCcnLqjgD68BzUfxfzM6fOxRNXjGmk0B9XQv
0pfnZChNgduVZNfZlm6gOgZFmTiHQEn7tuGAvaTx5BgUfnvQsl0sCGW8prnHNsQj
mbsvoGyUaD/u5WI0FH6T+8dgvylLQg8nj5XTcB3LCnvgK3GImG437vOJD+542Rkl
ka+iQjwapZztdjwftm40J9V+rbfgHk2PB8V2XNYH2T36bxeYFSywt0pjYtaIIADb
trXhe2OCBpvG9UUKBGiB03Ac+5onoHBcwx1DFseZGMwJ7I5lQZGrej9EknavQ5Ok
mSpQxs+VdxCge6OZyjWlZgOPFaKpW763Uq2Aq7imxr8i0bERA8GLGDHGb+u8WLBI
0CtzTIp7ZSW03b9b4BXJ8xEJ3jO8HebJkLtSMs6zR5ixG0F/w4csWnaIizNFMoK2
f6LisDn2IXC2O3umB0ZLTvhNFzPX1NgtSZk9I16JuVpmK+3eUUD1PM/xWZH6jS/b
PC46/8oFIzoaRfbdJfnu5pQnU3APcaRPfcOQldYwL64/2EQMoGKTVljjNoBLadx2
SfZ+S6QYJeOd8YR/lgfiuPP+JxCjaTobfCWiNIFFPC+dDRTt13kGw5yNloojLagP
KCdupQdtEvfR9CRGSfQudQktR7kYV9OZAoLmtkQsOrqHIQ6GMzIDVYbar43YfRqk
XdcL/3ItfIphxiSfUgQmb7qzcTrGCClMhA2es6txqhW5roS41twJglYPqfh3iuF/
XdfnE80HZvhScQe0ZPN82ck9XNBm5l2zdsY1sIgkul4w+qr+2cb23bicdyolnYqI
mQdDTU4jQqgOqTYeA5/qXeAorv7Zg9aJhu+Ndj2gUlrvpFmQ15RkyKfNRPGM8ljL
reSIom1umJmGREHV8WJzMYb/zs6GbKpq7OYVQUyMt7ltyQgsLSKHJg/KhwJu6YcC
lrSYvP3+bxbq58qcHj5AEsLjimVdwvuhQw7O4FVGH7cRQGyLzhm8OZ7pGNW3JJ9w
PFcIIeegoIjVSn00dxj4JVJDtmTSyhIPDNgQWnrWrMAVDd5dOq9hHma8zdu6vEIW
R/lwTkAUJJGDC5lkD9tCgrNnqSX7ZMijeO/JiCY6UvQ79QJJnmtKiRgSfptnt2Fg
ZckynA/cXgoSkIRhr/VtpknpF2uUQm5OID2bfmjUP4uJ/XltUcPYKSzSmsyawkxa
ius3W8eFcmNFYA4S1b8Va1Vf+Li4GPtFxUnZAhDlXZELmKB77alpJxq+MGPivxDB
miG8PU4zrw0c6YlFrZEVbgxOPSGjl7kYxw3QU/hAM8bM5iyQg+0ZYIBn7+MFIUi0
WFaaT8CV/Sby8quksLStKsN0Sx6yB4PWERBL/fLHQwlAPjCO556ndoGdOxbO8+Tq
43LyLr9ItrJZY154wO+yZCCXntJnkCMdmBz6HcgZjF9ngscj+4mex8lIFQDYMYHZ
KMjXn0K8ENQ9nynMVXWCIBAYp1gZKf0WuMoecg5bv6t2GR1AkMTa9xyNmep9vqiL
fXm2rgcdfStZZotjfvtVJHt/eORljNFmhzpJA/iOZ05mB9GFxPkqHoENGHetMMAJ
v/d8tk0Q8rx1d3THgbKYJT0T5e/pq5TOlsWO7rTkOLODI2RfbdVsJqLfz9nG3rE9
R/9jFC+FYhxOz1kCcfvjszc87i0q+kGrNpm5Dy5o0ErqGZBSAd+AJCXppYFx3rrI
V6mRMCEdfOmk4ghxhuvYXDCYO7b22Kj0qPwjEU7QqqCBfINzuEaYl7HH79tXamH9
MJkXICGxM4uP+YOG4+MFroD5K4ObM3iOCGFEf28q+mIs0SB9837ZSTEIsNdCzN3Q
Z+tsTTYpJDRS4/6KRFJ5EQAQvjwyj8JZZnnk8IUWGrivbkbIL9tz5K6hBk8rwu8X
Ss9mSIR3amc0Bg0/gYB3iB9pYGkvPD4QNA5XQzdzkAnzc48tUVZBB/gBiEU/ln1Q
G3eHOIjuTzXhX+0MqG90yVfzxIEBDm2U08Vp4WkIs0Uw9yu52GIAIQ5uV1j/9su/
svYdx8HIDnphU4oFl/ZGA90o7x1I703HQztpya45aUsVod9oFvDYiYtGgcUWHUYg
Zef2j50HjOWtL6OazGP+MnY9LNrpocD9cfG2suMx5eT8e495ABCqUmQGZfdPkzdA
bXyiSPblWJ8E1oqGrfetLjqOyRfhHPD0i32Ak5EYxEqHbziZ9w0EnPwzQ7uIDGdA
fdpc3zvVP0O3HgnQA/04NgN7veL1TpdB0TeeY9cJoNo8vQd+1/Hdi03lHf3EptPr
ZAiTOjxFCO6FY3gIFr0N0MV+AZWRxnl7kSq2sRWhDtlmssjOapscnTQMPFVCLLKA
fAdSKq5lhznwft9MJ6HYfCXNoBUARWIAnRXlFyo3wx2Utfe9mGijartegjjPfp+g
2DNiWocGaOHKRiNJJahEynauwYUAQ82BM0tkYrtgDZc94AieR+7qGQhTBs9fKUW0
ZUdUFbvTzkTQyTxp4j7RIAlx0jQ341T21bhvmb21/trCMAPISNJt8ZQ1A58iq3gc
AU2ZdIJKPQop1dKu/aM/Q3/LnWMPO/UdLSj1/LTpvQeLcCZfzAm29dZQxB+9GrGQ
XwftCJkjM83jimvIMka4ak39RgZwvy7IMUs+Q3ZVyIam11ooaJngZtGu27yKw8KV
C+YINQ+eQh4KAcdSmhvoGzUVfONIIvpIqfGwtFeA4cRRxKWf+8zA84exj9Ul3ozG
XrkEgn1QdfrSorhaAcW6wZhkHeUcF3nNcfEZxyP9GTQ7Ul6PYXzabXBm40Oq2tyT
bnXW48wiSIWzOh7OQ8G2xkRSx7wEa6wZqOJhQBKWA0yEYDQXpQCmccDZr5ECCaUp
/JsVDPPRosYVcQePUVR7ueVIyZZTqeThGIdtN5ebFkEEJdjRai8saWd5rYNjWJbR
AbVlBVIzRoGeBaE3HZJ+mhnrWhW8GB0qxLWHLqBX03IcaKN1vmcY7rnQ9/v3m//8
XIqMg/APXZNPW/YSo8BcRXQ9585nCTUi7p7EJ4i5vwVsRPDDm1j4ajqzcH3Dua8l
tn1MJW5L5GbPolVx2JPyJQeElkOBX/YfgBq+Hs6AV/MAG/RxXS+dMQCJSw4h7va+
JCBPKhL1yGVTBA3nRUBTWPVijebbT7X9m6w8LAQEMJa+FWbXsCpRyDvExeooF7Gh
I4ERYpyl8kJbQVEOds3tSLIFhBr1XBM2Y39bmLqFwWnj6xpCmghGeP0IvmAj/U9B
WHAMGtaA4O8Ugqp7+jKehEPJi5oZfe472mDDiFjRM0vuykYd7hFhVdrbA4jfp9Ep
ovfVnxILRtTDkMVLsw578s1LF8587vnxxVYqvly7DCHjstHofqnQVpTGaTRvXJTO
zF/uAWTGPYjU1opI9xqpsQxkGBRzfX7jEVFj0yY7jWRo3CB3AKPOERRsFTid+mwa
rbQFafSmf/3sOQ8MSRZXKdKep1dnmPZboFvDtCiZZg/yznmzeNTGF9DvuUUXD8QW
Bcki3BmpbZs1u9ELlwO/LOO9n0eceR0oXl7poGLEB6wPHspwl3TjMZJnEtTw/2O7
YtTFdvGvdVkaQW7CVjId5V5I0gUfe9rrddKwEF6ysm3QH7T06K2rvYCBg8ISbSNe
rrU1L7RBXpVWm5ikLTteKo9cqVG4qEBaiAdR+Iqo+hC8j5E+ToPBPSvqJPpMkv9W
REuwIZ4QeEx4gMVveyUeFZlqnVHspBUhgJcc5XL/BDLn8A6c0Xn9w9kebjon51wE
hSyzXxFg7sSTDIxkD81Bl6UvcQOK50FJLxh+ef9cWuSyUO8MdSQtxFMPtMdL07HI
MZ2Y6TFISjB59qo7MEsH0hGpz23hD73QfdcUp2IdZETDc+GOc+9ODpqEyBLrKxIH
pQTAUUBzZuRVAkRXMY4tB9/LgvQ36fLancFmuYvF4mF3dCTM6WVDUS80zNmqg/NU
AtlEcBLew2RLtRK6mUPS+Zy00jx0sj3FnMFIjA6GwJ0SGeg8PKxtTVwJAFU2yf5S
lsbzuXJP1HOg8uCqqIIU6OvriYCM0/26QJSPXmOf09er7yLvfEtA5/almQoisfwx
AasntiFeH55LVI+ffLwdNtNG+n2eMdnSkLtpa0PMJnewWS9r7roOPSL+Ilm84sdd
nalsPVzr4w91zMN97cF8/aDUD45GXy+oblfKgAov3cZfz+hrzEq+XUaP3Maa81jG
96XPz/Cyrc89Fz6kcElu3e28X40DsnIeRrQSyIAd8JDBGAHZ1Cu3vNa5JS6u8Qce
7KPYn3akxVhEJcwaiNRG0uiwrrskOfsDrLXGYTTFaXzQNZt4rWK/Cz4hjUkJ0Yc5
QNbcDWQAPKfyysNKDoqxqJQ5LtgGKxFK8On5uKvzURHWL8WHYf0cvMiLMil/lDxm
TXTOKD6Mo9pHwBYuExuFK3u+JHtyOOdiDnTPPAhurKKUHT54jfnl+TwsIeJIFhlG
pJckN03pjb/ljQb1MgzqokxFSq0mYo2UsoYwJcQ9AqQ6Tcyj0ajxR11602a4B56+
6ABCdLkoR7pOxfTwJ2M7TMzpoRsUEG3zioVXvU4t6UjqXgpS3pZSM2C6T87e2ld7
FgyoNCjDWfdEDvdJsra3k1ZJbeL/nPLvdo/YdX9jdU1hPga87tlH/e72VvM8sHRu
0jUxZdkyL9dSR4tqUBORXBOYeF1RHvUstUUWMSfGgvgreKfTqtD8R5q/p5q7xrqK
p5aNdEuP+ForY7WLTzTNdBH1a1Rv/nS8Feg3KeVTB1zZhCso+4tSM7vBc/s/iBGg
iSyiy+n7+3g7JFnj1fF2IiSAcl2bFaQZQLDWkjCx0AZJVnzyHw+OLDmMRX8AikqX
qm+iPYsGQpSiDeze0mWLI0EaTVwwiGrWMTnVPENXnFuTU+zBQSonxcLBu7DPwwa3
1iJm1YzDkK812p1Cp3WLIr6cw1zvqhUAWOj9PDTdMAL7iU/n+IahoydVgTlVqllT
GvdOqBmXFpMLxObWK2D1VN2VKNK5iIgDSH8odDCQ0gW0a5lWdFlDqt4BSHOGG9/F
7jq6sW2+Cflc8bFGOm5Y+iTFkFXNXjXpgoEqLZxovrFo65ZUQDawHG1xcNeRd8YD
/10KP6YARKhtnNFY0zGQnQfYN0XIcQ91Ztpvgp0zfuKMaCTiQVJkkWmNLCsRsRRa
t5Va4+MDBN5a4mJ0S2lqko5wS73wK2Qtrc639sVYCoLmaZEQwBSECvkiRAd6h7+e
5VhwhiR/RxVnoHpdsc3mFGd3dV90HBZFOYx9PMZKaHDwn7lTzQRZrEldPAg/nXj1
9bl3fdQ7SQh8eqkyuD2l2U1dWRUCkw3FmMA876KOgaVFwMLCF93XygzAbk/vSaRj
hQMeU3LlfomFBfWeNJnqAJ5BJ4fIHNDhWixv1r4oExmIGJJdVjyRTWVgbRmhUTOE
muRLtjrniqLnA8KpUOiLuRcWPF+FyCp6spW8oys4zrlRd7Y9vsQmhcKoE0hP8VWx
pJ4/RwRzrWj2UjWNzF+eWgo7AF5I4WzS5htLkUbOinxF6vQ2m/dexMivqg8b3j3U
vR0BsN+NuLwjeLKhqyknaAnT9pnVGKHmEsFHANe5zZ3rxVzC5Enn+sTZA9NIBdVV
X35uSDSyLA0J+sxLgBydJabgMTus3/Jpf0K51VPWB0jPr+bV+iuLtUMXNhd/jL/9
SAgkU+iF70g36tXHMbm7Ufbo8TVZ7Qmf4WRX6YmCIrbKh1cvtV3F1S6rjbkWn7nN
RXsmq05ATWbBBz+FS/TemeGzANTS/MosPMKXYhurbrD0NWV49+5+TNiD47vqcrNk
7jP8w3PB91ZoH9+fOSHUSYmmNLkHv/6eMbeO7h9qIcNP6RtD3abDQo/ENnmchF5x
dhs4qHEFafvDegntCasIskiYlTajgiKvfHsbl0dKbu9MQtLMCh/rI1XLuQR6E7cS
3S06JmPJA9wJGW0MOBHXJXMybqlnhaei/W+sbNr8sFuHR2ZRU72b1EE/PoTqgo9p
tCcIMdBciK+CtN84q0yVbTUlwpaSfOPxtDQUd1k0S21Bs0koufaGTxp9UG3zkFcT
6wIW0jdIMU519oo7XqHa9Cs4SSbl61aepK6AfY1vYSX0llXGa0cS7tAjax13e0pV
UMxBXmiayRPavyRLSADM+6fJjx08QzvstLrE9HIZUxxEaGxyAh+rigJb8DPh8RQN
PdQUELk8P2V9QxEKkAvgzS1epv5Qy4VYTGbO3jwltYe+wiuO3qphDeM32fnIyxop
5rYX9DDfHM9Pdw4jlEuLHlEfsILz1xRO3yCw/iwzCckZrS3gGEgFlIqAy7Bykq3/
HrSqwqkS7U5sCY/gsxWmPGIeghoJ7Fp8DQmP1avNO4P5JMrvUtEk1Pjj85OcAg72
goz44cynqabU04NVrgkDi0XRKjZ+H3VlrR2uXzHrwOkToiZshv+C+YvdpnDNw9+m
pC8w4eVbJcC97xDIHU2USm3+WwpRN1DqgIdLEFX1Dyg9Q603uFcbcDY7DXg6FjPb
n0b4cUYhS257cQl4U1nCcscCxCXDJIBIO207JewDvGUPWwaFTZi8iFSVlK7vkTEQ
UoPYyVYJr07exNi5spEMXXfdgWsf9hu4Hw6tL/1vTg2FwhtGlVfAqYPWchkJi06D
71IU5bXtArEUn5pfYHNojkbju6yqpLqrRoMuj91BZsxl0eFGie9RcbZXgAk5YU7p
rOiGxa/NqNzEB16BoiIg7GwEZqguJineKZ6PTDFgLj4u0PbndP1IUGZonU8p9K+F
0RUhfpcIAxPvxrhS03+Ym/wf4tCaYwtR0T9hSiOy4herv7OI/DDsNdZxj4gBItWd
e1FFK8iNeTzJfRxZ1xyuoH6wBIzK2SBY1cELry6l+oEsUKEiOwzhhIbj1SwJYXZw
c8kRNt6dj3Nmo5rwWHtMswoNrF3mk4oMhLayVYsj9q9/MrY6Ng81dB4kKv5Cl/Rs
RM++69gg8Y2iGfVZB9TH5NfnnfsXuSq1oNVxrkec1rcCR5A80igpAggjnR0hvjXO
Uc29dAezJ7BNHXqFpYb4EdE9YFQZNVVVNEmhhzCe/4yQmeBFVkMdD5atAB7gwclQ
P8O9+StUyUhY2PorIJw+UrJeAmKXdmBfp0Z0j7HTcjFBTvQCEMsfBSp+F09yF0Dt
4a0HLR/7vU+xTC5OUF6e6OThnyY3mKmCFeEP//v7fJQ0K0e9BMpiOl7nj9CbFio5
OvdOx+ksypNN94Lruu6iZVyHxh4qEFifjfIgjDUEUJkV4DVAiJtg4Yy/mULkRmd9
qvSFnguV9AxywkEpPJ87rLoSsVut+XWpBifHA02AxMtLpTPCrfUsaft7G2epRfNB
yGfkMf2I98wdmHd3MwcJVuvvMfmGPWxoQQfMw4Dx7A+z5MLzGdddbzkEj3+8NbJM
OVT3KGI1inQD1hvk2FqqpoomHswWlEWNRl8jr1lmqPGQ/6BXuM8/cYl/m1uPiddj
XcTvmvqYoYCKQZQzJkUfYdQNY9QBEuuKafIeI5wAQF39QZzaiGcqfGZX5BziofC+
jrF6BTmPT1zjEK6IoAKY/aL6riHl6ySR40+FpPZo//j5Gj9cYSUXn8m3N0LP93k2
rWSRRNnSjQ1k2xtJKh8tSwvwfNQqPKr2YqX0in5PNv2DgciRlX0EPYK9hJThJowx
KbVWCIlcpmx+bD453oIfit3sPQt3x89sL2aQF+sarWHo7feGH9hi8wM6uQqztm2L
XriVPaZI2t4li3jQl/Ewkaargpr1YpMbeeAXXH3B7M855DefdMKaxJqipNOw8Ngv
Rp93MCvoNDtpm2bZz7en84RmYZWXl2dA5CSSj4LqUm/8ZP8l55xx0/Hip981sQL8
62vG/PlDTwQGX+F8Q825UnrqiHZbddraW2Hhg+qSB741amvpIUpJj29Vgc0hpoEK
6iDPtBrDNEL7AUFn9+8rq3ktBA8I4d+L2Ocg7wzK/LOe/sYc+zn4QxblNkjilaB5
5hm72cD0aKQbwEkJmdwNA8NYdKm8WoiPDMR0mVxSYaSeIJ6XP5FWhrqGFXpAWzYe
p9TOJUWITXH/HdGYnS2Pr3pj89dJiReQjLpwnafAj+wnMvTBL35hReQOnsBc/PcF
LF/yoyPPWYPb+WxbUCbxJgg7+OYdT+XvF1o7UpG/SG+fExTu28YiiI7WD+E9qG7k
lSURoEX19gew9jML9IO2nrhVgmJNXQQE862DzEPUYH2B/h/1qh+2Owe4vHhw66QS
IrPr7/azhaPLEUwNBtcRQFru3oNrA0Dpv4taqs9d9ZbrXfq5bjkfNlBr6FZE1aWf
ssMoLXtlPsIDAs6eMpsLSeDEGzhNcvA1VtnlA40wB3su7BOdA5K7kvy5um5madct
aiiDiQJNIYOheNKqr5UcJC0ikyTC82L+9gxOiM+LXH1WwHAbyUgL9H5SAn5qwS5J
3u83QyZWQXervbR97qQ/whS7zeLqOrdOnH0tmSBAuT2LrFmwSK5WFIc1GICQjLcI
F6vDrW23C+KfVQKDhktf93f7Tex1TQN2uL+5mfOKNQQu2EPoNzMvjFg3GnvFrUGk
kJ98hE1LGOVg8OhjPQ46WiMjyem698zPf0BUy6d4xVuh8dNuljjc3bYmiZeOb/76
RAUTD3AuGBpQTSHy4qSGLYKysuxVO3FsDgUFqaNr6MMi+DdqqpVGbb5kYw8c9mBY
uaDyLzb6oGLUMJvuQEdwVPCY2Hd9XelRM9upSm2W7VahTtFRu6V05wyis/RObEDo
T/tOlbeW4D3NU16iN5hZVPOQCvIG8Vl4NtzD1sh9r6uiKEcJn6S2KiQYsqD+/C2w
74q7vjZH4KJZTHAd6cw9p4iFDJHiFGJSVJYkzF2eoaYU+O6rPsMqvA1+li+W2w0b
CbZolc62i4IcW2EynzzrxKJvGgdvFMah7gpEh30NXcxszkFreWDT488jSDRQR2oT
SpZO4PANzKDvBwflcZD60FLcuv5NBalB6XtGBn7mNkH4uXWWROpr9ok1IpRJ2HpU
r0xXwAkVRB5yYYXEuNj78e2eU3tooN09KXw9iMkgFgAlkTEwiChH16r4cU2TuI4Y
kq3b1M//EsK1BDBywUTMRo+3nkycwS4FEPwuENW+twyz4yJ82OAabQxHAzgNjujs
KEINepZW6G8XA6V5uW08TGI5dR56AbB+K/Wwzhu45qt6TYsz0A1qGU8mq/bmtyOt
DcH8WJXoAJLoVa+iVDzdHHGZ5HXGP5VNwb8lv21tr1W11SYDuYXQaAjtyNXlecf4
3dT9/J/nAWiu6414fpGjVlzVFBjojv/YwBlyiT9RqkcMbypyWjo9sdLAeT3Z/yNC
UxJSY3HRwtysHHbGQVmuP4zVicKkoea8v8+QscvLsFlS+CbkxKitLxXeseFy8T4m
Vrck5Zq4s4iRsIges4UVHfot4z9vscbOJIhmuOgZ2ENHxGOPaAFQ4Q1/KxofmYuv
eJQlqZPZlqbS+9BB+H920DyO5rPp5GYCqg4+BdZW8TYDxT38PVoGr4tyFz98Ucrt
Ro+2o0uZQ41FHGRONUXgocpSJmasDM9AXy8ybdXGAnBPE9Vmo18IuKDOwuY6Uk74
eoedLFoEpJ3td7RnwYYup2Cof5EUUPcgZkSKdDIzwc+ljxpfDz/5/urTzaw5Ifts
sSEibBOywLl8jHPDj9NnxAEYD1yAWy6Onu1DCYyznacHwiFKTD/jr0Dajb+4A+ig
SH0lFNAvgzUdTPDQTNQJfmt98GYzg4lJYnph16Q8HyA7ZgWORiHzGIuPNOsYzNQ0
nIxKpLR2IoUIMNvUjwXAsqP0eGB9VyZKz8uHtim8jjxnTHvHzCXqRzYIipji3oIp
HXJUav3QfYjkynuLE8SOBBnEGpP1M5a1uZ8Dnu2AsrJayaPK4Xt4LlD5qwjnOzEw
mMU/w+VkPfsfQXwVSiv6iW4bnrxhLgMxI8CtA7Z2YZG3n3zYhKxV0z/JP3hHOkiq
L90Itn0DODqDaL0+oBc6ZMd1/irL1s6Z9653FAwPVcIP8ZeKsxSK7X29gsaOqxTB
N4GHQkpvYl5hnroxP5GbA4P7SBtuSyMzki89zjQO5ZXa+qCN0j4+oI8Vrv7qfxqQ
Ngem7iwuMasHpqg2OvRstDZUVwLSoYf/Lqr88MA2slzOfJ9kqKEI6fSY16AuCXjU
j/UiRUVG0DF2+JzzlV0dVGvQPTFgoVwjmyYEYMs8VwbwAdYvYPXIPs7fNfeftLxH
SeRf/Ve693T7kDsORecWmUyF95qzxTbL9OxVwd/6m8Jyc8qI/g+5st/aKI4nlje5
dbdzVhM7AFolqTjQfVRN1LPyNMPDfjElXb1VvYpr5P9Vh0okMB5YzoDzBS8loTVL
ezlJ0qIocfxLGGztkbCrTFlSw68LQFuGRFJod4laVJTXdKE4zCcFO9rZzFExb24F
nHzjCeQ47kH7zEqpWG+rh5N2+qR8hzp00oUsJeqYrtSgsjz5exurppoE5f8KtM8v
rYajDKai6FEsdWsz0qAFBN41TVOg6IO/CA6Lz6OAelajyV+yJ3xB8JXaU5jB2vzQ
6zpKPGM66WwT/9BWKs2lPmB1Y2tOaQAwH2mY6emJgtVrLvVTxpMw33as3RsQs7sR
e9cO1/N4zQI5682P+GQyFfwl08mWjl1RNKttGxIL6MhV3tMcwbkGNO+TbxkeD0nf
whMm+gClQfVwTYgCBb/Sio6/rIkyVfeP5DuVlhNoH6EDMXpQvGEOcEw1PcvUkKwe
oXVaEYQ0HHrIijTBVz064YJwKzbJxqquD171N46bJ8jd54h63S7z9Ed2M3PztJsU
k2F7+UJ6cf2RJFry/OwLkTCQY995fFxT87TFAI4C7quE+EAS7dKpb/qRFlV8oRUa
hTVoAOEdnNoAsdazde+GSSmZxg4NrW+twyoiVQJTgQLXRyM3PiW5ddxNImwXS3MD
AJHsd0V1nns3jwxRUAZtDkNvkbaDZnNd9VWmILOibeV/UM/sCrgBKC/eBhFdPRLX
jnxQwj7yAX6HYuOitkG22t55czV7D4VboA7hEFUbrRDQrdQrPHAEnbyRPQA0DRME
qHY1jE3QKryQbQLE/nxboBvEFBLKu9uzEfDNKAB6QaPqlQAa38u9gakqUKTvKIpc
vNJcS8FPsVoNEjBTcNEDxV+1wlt9KBIKJEUm6O768WAF1tUiU8YJ/jNn1jj1Nf6e
XXBpK2WHZrix4heZHLbqBUg0QBBGowjWk2IFPqaTivnr9QXmx2jWoFVy2BsOKZ22
mdY/VVXVkDEyiqJVwnVxRKGVYTdwAl5IBmd1yBezTIpwjKteviLE1AGL61DqiSqv
iF1kMIrfbJyq/mqUB8j/rV1AORXUdAK+aT3vovmzhvaKKwU1+yX88UQyBQi95lRt
NYqOwKdn3SVlu7v6EEZumvIVmyr7abpGjfaQ3FIxEZmUReUyCc1ABeSrQz/suQ5+
Be8aiqMYwN6N6mo29bjG1dh53ApoTgluwkz0ZSzFCcJSjOLw6CviGXRmEu6ZQSGI
/yAUjFeQN8Lhwvvs5uD9NtygqRcEBwCd9QhzxVyoF9Ah1V/O3TExLUMOhMXxAzCc
Qbbb0+DRR5X1CeruetiOg5j6qk2ijS8r+zZN61fHpFG8mgzn8a+dCWhb6KLBj99H
zJBXOoiurDUv+7IwO5PJUc7c2cC/QhETfyHLWIQZZnpoTPaxYXipmVEZ0Sm6q1Ww
hA4kDRwOollL80C6KiTqAjyXafKvsdfBvPgNA/K3vECpF5UM6AOVeZ29Zzhnotzf
g8+YwvPfTA46PKBogRzPV45nRzQ9vgiLhAGFe2JiKwpFENBEDBEwGkl/tM0lz54c
C4AwoRXOuLj//9Si3EAnaNa7HOJ3kLDSONY2omZJDVMO2GmYUt5ozvAgoxTkp9Jq
x9c5wOFtRX0JfDy2PjLiucbzIYykYF4tmLucKRfOxBXNZhogabCiaXol2nxnL4nY
AhGddY9dVCOpyXt0n25bGwcizX6+EL02+81YTb5Vma4hnTgbrGfVkVGPc9oN5eSg
6vVXcl42NI0oKb41wEMUNDuE6JuFs1lcuusEuPa1AuLb4CsvxT+OQNpnQXVDy9NN
vu7k7K6gx9JcwPEPLqOleMIpKz7CmbVgMG4kEJIDv3ZA7/ZEoSwiJvktoJEhnOz4
WTYKaI2qbIEK7JgE79aWktlQrZzPQv2FdCXPwKTkzmgQcy9JWpyciZMMrlbtg0UV
KRH9f3/jd/T++ovbZv/Ic9whAFCad2c39vKro5ehPa8xCyUpTjgjj5xmc18fiFNv
5qohqtVKtdSCHWaQYG6VF2/WfemfkdHsHY3KpgNhWX7ih+7r2oYcEms+FsHQCrQ8
37zApz9XNjvAAXqD1VZCNF7+vIPoi9rfXUkoPCo+LXMj3tr6jZ8H6cTuQyldkEYr
uQak4xnSAmCUi5q2zbIrkTKvlP8Ug7BBatx6tfvak8/Yet4KBJ++6V8FwjmB0nck
rmVWSLA2koMkxO4dxwQwo8V3LX4l0l8qGQSTmKpuDH+x2zKTGYGZ8RdgReuiZcrr
vp8IhtIWpttnxcCLQrsMYT+QDf71I69XOhxO5xi4yDUm/1wShdJTuMkp19HVmc+S
WT0Bg7/7r/20jgzkYvBHwmnmuXOsR2TE7AM2sZlP3Z8BTKihQTMiwPbF7kIDgEy2
ZAt1DqmlGCG/DIjyMh/oJuUKb/Ovzk9oK5jE03G8K3ZNUzP/qc7dxsf8lpt4cnNA
dtVMOgHxxLpTRFckerLgBSmfAXfue6j5Squ5tZQsTJp7FNn+VgUt0lRraJabCe8n
a51DsRFZmpEqv8tTU3hqEbdWE9uXa42Ku0FpmZMzMB3+Nwa6pi0b+kmN9lF7nhy8
YEG/214XkpTaDleo+ULDqZzySh4dyfzzd7VVmcaylIPZ7RUwbCUCfOxTGAOjIIkx
JwoTolP09fznxMT7MsOaYbxRdGuA44SLzxNVMyM0A3riURGEddpxVmj8XbaO0JtC
m1n3HZLeTR+lgAdbt/Cnf51rBX2jZA/E1FTRuH3NHNC3QWTo9yva3uzT+cYbyfzT
aKYsK/CHw0ttxpAp3/yKeTdoruWO42YbwkwVY480Wk6BhVfNp2M+uz3e+z50tgds
8fnm3i5Vt03loys6MNTJ+0GIUmjAFf+z9Ph3z4IBVfFpKKVZLy3gXKQm66hyDyaT
OHDYY2kdjy4XBwk9f6vrh6f7io//9uoWz8L5f/E91WV/QCOn/Lez9QeYhMohLMoY
7c9i8c4IEE4Spf4LAfO7xt2RRU3xGoq5MF7kRGJS81OpiDBnG5p7A8Hx10GMVskI
EIKHyPt4CYJTjuZ2A5J2eLA28q+qvgoVhsEEqqYmXj7IoIBVLbCbDa/CpT6vlT7f
JsgvGClYZGeauagkrDbtv5LkROcuvpx5TIo9IzZiGDG2Ua1Bca1i8Xc0aT+NX9Bp
FWJRxHJ8JCotXraZc+zUq/8faz8dCZLgJqG7XxTHt5n7xKmrb0rkCO4dvf0Uihgw
k7J0juS7EOZF3MbtPvVrO0QahwCO3Xnx73ervkN7PIVxWAaBD7+a+BXPJvT6U+Ph
26VaMVQDbiq0GebnTK9lfSPBGoV7xG6SWunKuJ8lGeV5j0eCSKYSIY2gYvaZ2DSD
hAVgL+//5Q6ZxXicReFdQYYIBb8S/Tn2cS0CmJEbxHwJbWFtojfvciolhB+kkElY
LVaGbxjDKK5lgT+Jt0FStvHhrqo6wMnbAeUWTUj6c97YHd+i+qnxwKLIbx6St0tU
bQcYjlQ69yQzw4Nvme2NCCcXDNX5zaxgt7rp9BtAK+iNc27FEfinYn13uiHr4j00
tZDx1qDhsLFBuMHF+SburWBQnpORSLGRjBHV9gzSYCOKurl1gMZnrEl5MCjaOuMn
66UwgqFtOJgAQuF/G/ibsJDBojyhPKQl2quTC6aFB6bdOyPPGDR1NRxzEWcmIWs0
xJEubVIjDvt9p1hUUqUf4FlGKA2ujlY46+5aLbKd5Gtg4SJ2WfSassn3t1UKzOVy
D/x3E8kwfpvh8/TSMMKadJNUIfNhJAHabxkoZcskjHTaPKN4OraSWjbgyIS/sP1i
xRaJ7mZt9FJOZhqTh8ep70Br7M3Cp/OsIB1V8LajZQZVYUMl7XjGzcIFRSX0inEi
jBsJDOTd6PEVoORLd6I09hSBrlzyErC27SFnpFX/yNG9OPgOebjl6whVRRgMNjDb
xEvE+LJ2R/n6r7F6qNoATCdj78EyOx0GG04lgDYsYxpvfz1MWb3yR/ONgsPCDffb
zfZOXDjIBy7ieFjX/AeHXkTHFt2Uh83lXYFQffOdrqzb/kU6qhyajLj8qGDQb8wA
kDgc067ZErFlga421E00KmSz9VCEc0WjvpU47dno9+9uZkB5KocBEoipBKv9kxop
McAUUAdRa3nup8PYy6thdsUkntgfOJhyDtWeO0AE3Hv4rKEngYsQVwCRd361ehZY
eHrzy6mKVCEo+hvVPfLvPBnBWGRM4MI8GlfWzVPqIE0O/57YIa2tG9Pjh00FCBPz
utg7yAQd0GQnzhm9iItfF13GKGlJHtyR5gOtq4oR0IrQsSSzl1BMFCm8WY2RDzuS
3tdgG2fPsGOUx3XKu7R5D/KaoY2m8rdujSgvcIix2JaWmHTGA9ntP0D+D1uJYxTy
aTk97wqe0dGPkStJkCNu0dFexU7W3q2/dHoUy7tBH9Yd72Hhf/PgwXNxh8tgc1GC
QS2OJLRS3e7s5sCRxGylDL6hzxK2JDBVYynV2WQtAYH1CkKZ++Lfk52zgSRPWwXc
17IoAHFj0BBV9+7JUAWHUi/v59cZZEYGL5e9e8yb9pgYAmlAk3SGnTgB530WZIVl
aQUjTAZ3cLTQ5XLTn3i5aWZDzUCv+lC5CTFCc0QSmwOJQ5Iwh0n6CmFL8MSF5YcK
kCTPGdFOCIzXNDjmO5NTffwFLT/O6DU+ZYBgDa6sEJFUskcOjlFTOSrN7+VbGXbc
3RMNRisxpz1Wpigh1JFqAVFyPhQLh+vbf304+azZPYeU+E31NNXN67kkCDHRJHev
m0lyDWJWi4Uha6Az5CDDvaJFmxei3reHSgDs01iPc0LbextP4/fyvLT1zcEHK+N2
nDXTgB059eq3+LlvVRP47aekOiPIUoa6Gad48OGX5hW7MEX+tWvayEk6uTfawwrs
uHhE9uZBMphu8MRhj+YLB5ZbxudWa+yAafeSogW/+1s82yhs9k+NPPSdB79iScER
erh2JCZdh/+TItZAGBZXTD4+pPi2GzCtXliSgLeRxRwnIfmk8zJbImroHceec4Ww
1E+x8cbGf0HJnFKD13Rcbs4HBJr/SUxaD13SyVPP5FoUzM2/H2qEUa3WOt+AgRd5
3wvr8h0OVhWrsCymPwDSJ6qvI8RqMYtWnwOUGOwC/XbrfVpJpDUH0not1oQPDsCC
hI0mmz9LvtzcwcbpxHhfWyU+jyeGSnY9CHuJJDkC4A0pDj2lE1WAyiyA9pIA8yOy
mjvgDE0yG54tAU0PaKtgoGaDNsewGPieDS9SVlUUGQwGQNKevflsl2J08hi7nMT6
YbkZ08wAtSJx+Y2roIIWvXlO9epg+i/Bi44Xhp3lUscdT9xR3QlyKQJiuiI+VZl/
M/emspFh2Z6YaM3YG9tKw3MDwvtH+cDVWV7H3SWF3oJYfw0BjlSakuwMGtQTXbAm
Fu9la3Wi5pth0I8EHI/aUGhdWfTRH6zA7HsHMPsLeQez8bk+VqrRyT4ILym1qeui
9iFkptpGjhO46IJ1pvQuzshduLGXXKj7NWzoAF/bTZPaPHcNjKwPsc/0L83bHiQV
Fr/cF5Xgbp8fnSw9YkfvEYTJ/TU3CJkAtKEt2/faMIDiydiBqnDMvWwm7e/Uc1S8
Y1hX3465dvtdSNcfVJzrYtFshIz8rhxMUsP/hJ8OUTF7iitTspRWg6aUtcbJ4onc
It/TXF4HkcFq7JsqIaCNjNol5LHGoWKO+q788RogEfcrqzoxAa/Tg/C+8JPE2Ey4
PsJ2Zd3imviVhcGc3ZuuLXLhdfECKyVNREgfZbARKc0zXR88cKtRXk3ITrITfZS2
kfQzzUkItCvFBxGCfyB6+pgOA+Gs44N06L8qYmQ/zVNWColaHkK2IVHeVYXOR69u
Q63Llo0GO0wzTjpNezpA/gp5DJ0nJRS4e1lOYdwCMQY414kq0xBJdXfWvJyKQaFq
yBDocolFUrczTwOKnLJYH26ybolbPTZNUbTdsKDeHBYzg20j0o3c6OijOo17wq3D
7E2qHzlD9D0hBkUGoXzlmwyo1onnCAZdAG3OorQ9PDEOpayaSVayw5ZTj8MRBtZz
UTFIJI/IveS9Qz31sIJN8QEeN75WEdU6Vd3mDnTPhsFBIIVexv2UteBlCgT5uRn3
oxdn6bU2TFFT5dLTzRFKo52O9pgpvz3bnxJYXQN6WKri9ubS3lWunBp/1ddETa96
1XuyNdk9kpK7rp/Rst7Nek1WaSCiD+wb1pdLIWcwd2p1QC0SmTULx3nzIJCA/SAq
ngMF1B4LVFWbZu02rSmcqiqLmReApFEkDwb/K8R6ztS5pVDFcpI9nsT+ZwGGRHJe
8jqqKs54eQ5dAILy03bc8N0E7GqErSbwOn+mO+zOjAmHaPt+zvazWZtUDQnHVHqz
Wt7fSnxiBvSrp9VWTp9Kom+szoph3HJbvTMqnUsZyNcBAlF0CWlajG1Y/BNlW7S0
zwwhS+WkyZj1SJaz+vazqiIrLYieVjRszrxod/9/7yRiEcqM4JA7rRHjfB0bChrp
3WNVdFnTJVll3F5iYjMgPMSQ6FE7jgGbxiMmQ/IK6f35BeIgy2IJtkkQ+oD1qf+B
fon9NnYWzpVtY7eppSVN2T5k587gf9cJB/pceE9mTVK4J7PuB6nKHNkJ1nnu4GT/
rqOezaV1rN/71ZoknsZOcOw8pJ0R+Hg8KZg/wutp9V5iNWe5giKMj3OnEyDCOZtK
+tWrmBAIa76ObT3AmmcdEKLLqDcQWNqrMUJfOKD303xPpz++UHuP9qRq22z7mpR/
Vomp5onUMnNsdZIpO3CBY8nGA/ltCSQLFqqtb1syP83kYVIjEVkGHM/rb6EsH1xk
TiVxVbL1RYfkPulNTmt+MTvgmiLcOMJVRB2bqXhtL3kcEoD6+EufU/0H4WsVABH/
eSVs+jZqBwjZZNOZ31jPrzOOK5uW+HOnLXff9Uoani+MYiXxUp7BuzfJ8eBDv/Za
+g+XZafGyRKcXuPz1cMAhlVTa0GsS8UcZkVxIGADpr9ZuVnOgYp4TkaCWJmSI0vE
SAXZmT5YCxlKZM2IdxmvEG/G4SK2Jbw3rG+RVY7PAkOlxEh2FKvbKIoq12r3RG4p
OjtDUtjn93A3rkWE5z9yiQhl2Z+RJbsd5dopVkPOO7cVcO/eIF05nH+y9xDJY7vN
YbdHHmBnU1p6tHBBclBJfBBNT0p2vQuEgPeflwl4JEK8MulFrgkwFFDQkzKyeXDT
MXT1dntdigdHvC5qzNtt+a7WJ1rGURsbgVOgEVoijGuqcHs8/fbPY47Fw4FgQHpr
6Wsygj1robgaSU7LQ7r90t7sd2HEZdjPl94oiPxsI73BMGsTfGNulAQXZU+EJL0p
UD72cnxklsndRnpBot+Zore4qDGJvRkZlWHeJHc5jY19SEHifBNyQQvl2I37tW4C
TsEUrsNr2tSaEW4Y0Tz0bkxO9ok8mtWaVIny02T82LBscKHH4ADIiB5xbp6rHy6i
q1/NCeDg1SRORl+3BseRL5LFhbYezl5HtwZgFv4cDKiWIx4f3WefOfPVhl1zU62/
wMsrWfgOz47+32veQSvF3A9uwHeFHwEE0Al4YzwqymwHUBMzvFUIKB1sXO/QwGCG
JeK5WWEbU7PcR8U40yIr6FoiVCpNv6t/0TgAmpcIAlF+WeFYqT2yYzo584dNvmlo
GFuqnEcGbYzAAIM7bvtwK+qldrdZXTT7qBpu9ruhOmza6R2KSTu0peRBxI7M6hUz
mGY9CJQJXnxqwKFxGSUmCUgEfI6AlU9Yi7xGV4TLAGYgTzc2hE2VD3TGorWG8CVx
0fokA/M0tIudHzH9ckwe0uwIq932slKbZhN/hglj05KdYqylvbqbdhYIeuLvTONB
xThLyFxJ3AwDuM73nRUlLioxIA+X6JhbeOR62451myizEVdH/O7awu4Ji4/S7Hh2
/mfs5rr0la020lJ8hrqjaPhUVhjG6Y/0+lsVy1MefdaYjuLrljqrtIcPcowe+uNf
TwOrFwN8ZUQ34xenN7p5dB+McRXJZYF+Mv3hYKBXQZgJVMD+FPMj89kfGseVv98b
MECyQXLCaTuDpAw1OnKvTqEbyArUJYiHVf37cBVxf1yUsN0/aMTzxSx5GgdRZPZ0
CBk823TC4591edjj/eDJlhapUcY1Aq0saPqRa0qkQFvGMzYX6CP/pdB3FH45ENmF
IopOVlYpc7Yd+WPvAEW1xSVCg632TeLK41Jz4nlOAKQW18dR4qMwhp6da/TETq10
hGPVL1/nZNKTzixWlHikT1wE5FemHrNW50BLISQe5XEKdV7pVKfSbjaaX9S8nbqa
AEIkTU2RIgKw1ErzO9air4/5gk17CDmK3A+gvhd8oUKvPbpzJ3uifrJY6zwFvZel
m8TaZga/nAeXhAH4xUpJeror6fQUqEbmpvnR9hU6p/G1nGQXIYN8rb4gJM4xKWuf
tINRKfgDxgI0L4J+tBquVHkEdEdG/2gr9Xc59ESUYg7CJ9y/O/M9hOhgbouhL/9G
HrlnyDa9RkE006mCAort8fSpw+bN06/I1JBAMUcpZ1tNGeLbP+PMU4SgVM5rbh3x
khP8zdaQEnIVP1cPTJewDpptty+z31zf4yqp2Xi+PVszBV2vfbCC8LuEe5YxwWQp
BHvd2CTnkYKg9ISWWjnaDI+zYHoTVwZYy3MTRXMsMkyK8siMljNb/H2fpgtc5C4A
1s5BCVgg8BLoFYU51OQ9dlv3H7iaLdK0vgOiJZR/jUrCfvxj6gMlhoVUKKVokVss
1atbPgS7SLFk9reKGp4IJgUcsR8cpgqVuw567ahAHpDHgnBkWHyhQGHcuJTD1cuq
dj+BklVBwu3pRy0ez7G0+OyQYkdsE2gOo9eLGcKy/OZgirtc/b5WFuq77HQ920gp
5OJRPuFwQsMnpqCgiNqdL+3FbA7pu+AxLPqhFg6mg1WCYebqZfchP45yfqscKn2y
rCtIs1oBeVNDly5cw3ytw0J2JV6HBZul2VrKl08va+8Jlpf+Th31jnPEFzyupFJS
0MA3Dkfh3hTM8YJUAcVh7v6+oC4GmwZnfOWAjIs19TQ5QoB0KMLlD2bqbiEf1qGr
AL+cPoQd/wUoimW6kbrvsBFYAN0YonqqqTIrpP6xz6h7Yh2u0lPTNgrqdpk5mmJN
GYuqDOWK1n13FWILyHnc4Zax0hOQ6rmwToiS4E5PN1R0+hLHin9ywwzuZ1mGxqXb
hqvQTM+XukOwop95EG4tnaEGXUiaLXJBIP7xceNkaIXbauKUnYEGCr6vjLJmRo7W
2OACmC3wAi8UR3P3IZeoC4etZaaeKX6ZcW7eHoZoL3Xo876naisHoIz81dKcxuqz
kMjtGsAknl5Kk1FSLYUK3S8ANjslsKP2Y3aDxklnGTIlT//NbZi3BaYBdWJwadGK
v7ks8MvQyaR2qPbxIv1tFp3KMzyk4MmAaGKNTTcPXWgbh+THI3ANWuyFC/7CXdtl
Ht/dyzvhT9ScSnPeyAbw9JdmGVBgtgkIOUsayR649EA6o/6HkzjmjQvoCzerT2af
Plusmp9PNkZA8IfBLOz9RvQZAadfAdybQxhyHeNZwj+3yi8AwK1OpoPSqRQ1NSl8
QkHdEMyqzRD5ZiYvVrxI7th6tWils6hlYUfc146DIX5AVd81fR8cgnfDpdbsOady
voLi2pynMXd0St8AUetpxAanC0/VIRhzyXWhTl/6dWkLCsgtPVv6K+C4evZ0N+ZX
Yjq2RgmjAhg0uf1mFJAXwZrY6ql5MJu5KGm3O+244zfblQQO/gGMg59cCKCkQPVq
P8B0tDNDII1h302Nbdox/ahuDGmL71TrUxydcrD4PCmo+XZBGiSM39A0exZvoaKf
YiUIv/V6XCu3M2S+sOdBXCK1LVZMl3/+/s4nRFEklFeFhbM06ZAS7hcE+o5t683O
W5Nx0/92QCkKm3CMCpSe6qzu1a5hZjR83pEi6OakplX9KGLBkiFLwCDDrTvIhVfC
g8rXJ2hm6YwHx9b/0KdBKB+ovP6p/VpTzrVoJJhv5pLqsk2hobVep9KGVlg18v1k
Nb9jAsQrJ5aYaRsDzkPoB4FVdmakDt05DtrXodZBr12sj9kNEqPM4/TaVrHLYpYT
4EMPh9tkIi5kZufffmwaQIRzckonBWENjP79QU8Aw9Whg8VAZX8hkf0qW6clob8b
ImQtHsc1I0ENH1EN9Jbp7EJiLafbc/T2SEH2Wme8JHgoLoEeujiCDBI70DmItiH8
73HkacL8giFUIT36+rx5Rz2fLdjW2QUc6eZnFIge6TQish3SPekgrJI20U/jtL8A
FQCP2sFAV39Fg7hoeqvpepuNtzYxCHmW6vGy3TZ16KoP3ZTRilbJPU4eMAyiNqus
AxB//4T4d7jYIoxZQAbszYvjUkaKMqhyH9aHS2wZ0/dIQLWeRop88EgHT9OtZoKL
dqTDRxelTozf7fa6t0YslG9uqfsOscPTBQRwgsPa2hZdsGCwJiJ+niAYLute8PIf
ZUId1Xk5JFP9zDFNlNQ8ECHvttdcQr/dCAFdx+ILi8W3C0OlHGP9yrH112CDDLIJ
cp6r/vvKD5qTtaik5LN6zEtQE32Dl4/SNsZ4kMgoYTfXUHeCpsS/dWEVUna7wwXK
ypzrRcd/aMc2j33Mh7TRLswjx47/xY5TyJBeIJMt0KrgCgmIyO2yScR5ILpbatFb
m6Br/CExrVg9Op1qiaCNC0JP1kVyV+o2vjqO2hnVPTHGy3vz6dcQ3WZotfcKMTfM
JaAHMQxcRwZQFXbqzvpCS/PwBypjI25UG3ei9XKBqO5H1wKUQL7HArRS1hexcPl1
QAHbLTD7f/8IuzFYGLbCIJipJaD5oW8Xodz701yFUmRaHONJWeadxeZ2toYALeco
35DPl+a5rNO1cw/ovXcZNLkkq+dJfJp+eCYX367ulTVY2PfAOUih9xVQw/6RidnC
2Xpq4Rxe8ZbJgzvS1MzvVQIe7AvMKpXu9PQi3YSTyuSHmLRbdNTptIFVuCavYlT5
EIlsAp/8rUXdK5GQp+V4+x63uh4UhtHw5RQPOSJ8x7eUXiSiCeiKb4YOyAnQZgz1
ZZTtl4zWR2qConFfjuId1MsR84uMHtsG0HjjCpjm/DgFVASoeK/jKU8nDWrGN58s
AgFl0IX3JSAlPUarqJ2v8vfFT6BAlQMCF1aAdRzDrhN207YxAa+4x4KSH5j/FHpG
Ue1LQERJ6q/r9kk7AmBz8Sr8g8e8Br2On/L0PHtbQpdCSrwjM+7SuG0euMqpuldD
jkKk4xdzquLyxtXW8sEovcW8vI8CQxxJbqo64HmgfzloHiAbKNursL0WJcrxIGrD
Ro+HBYrVPMhYCg8p5D9MBRSuR814Br67YEWJf+uxth1R8egKW+8+bvChDcLhpswg
1c1iNzz/5EI8Mu4Y6Iep/7adRvR1wyl9am+ZjHB2STyubJu+NVBOopoccwH/YryP
V8cOryTmddz339Xfh8k7+ctg56SKQzfZITQAT4A8T6LlVytIwTLw61jisgi8nVSJ
DnD6skW803Vis7M3jtv2RjoEh3O63HlX5LPfz+Ym6ts4O+XEuFOvjxfsDM0eLGf8
VccRro037rh0h1AEDTUQryYMAqhOMP64jIAinysCitUKldBtPenMn8Qbt98H4Lva
skaKTfJviWbmXrniS/IwZfNRz6gNUiUX9oybZcBsq1eWbNkQ7PxgkSlAuGCh8pDj
pWVnW0+3Z2IP4rh74qcMBWS7E5A+W405vekf9lrWRe9SPeh/FILw6pxpQuoP74kd
lubBVUHrLuKeexrv1AckS/zGGD3/bpBWRgw1ihwKt9/6kaboWo1H0X57jbKukk3I
MI9wTm42eCz7puDwe8EPxBA37gFU9GzcM3EXuipDMxdZ98AAQVDaqMElVBsIQqIG
eGeInMf2euSvWJ1saMMUHtrV7Vw9cDflhGZejxRmdtsVycwvL3iLe/dL3MN10aSL
weSsENKFMyJ5YgflxydUg02GwDNELyNY5W+yt6nVVJ1aLqiIwmx43nL2ak4mE3y3
ufmsS8eL4qOcy0PiGd0VAE2cnOIDPrCjmt+9FBiw9UtlUx5X9pxN20wjueMFaFHP
5GM7YuefPTrOLb2pnucbMjj7mZZWc6EfXClcQACDpevvEEJppxeiwU+IWIjdPGSr
z/HSsX182Edo7JYznB4JzgItZt8IsLtwMk0r9w+TLgIh17HbW2Pe9wxialx6Xi5x
xSPDTfdFyaYz4BsI8iZIMjF/qb15GKQhHsXxJmeY0DZAtonHyfQ8CSPti2H1hgAr
m1+izNU4uFv/2wd1urq+kzGaBE03hhWuTngsuGL6SqSgPS9b2eqeqmXQkQT9+CdB
8VkFi7G42kuQqmUU11D29LwcXc3YVn9vUYjK8yQyv3msBvYn6uYpp2lJOzSFiAty
Ntw/29/fktApT65XT31XZCBMEzAJOT691+IsguiiQfWgcVdH1kaF8dIYYGIR1JjL
mxkuTpcfHhgpi7HlRqnECzsNODXdq5uyAZatied8mP+DSilY+uFDd7mHt3/pf3os
ad9xxeDXoimT6pMPNLzoy28W/t11bduFtlKJXR+T/p3vMW65AmNFZeH+fGkm08RH
thAWt2jE/HdgcXhFQiwqlb/qh8FZXsH5kGIipqGcy6tSmDx569ub+upHeL3xnkYX
DL28ymXGDckmdFQTdXzm0cNECIhs2pbgEB2/YYiFTqvrrf0Khs0FXBMOLwO1smGk
M4/aFz+iCR2yciYR8aJnx/yw33KKz4pmsVh/68mkAzrEB/Y7kjRh4EZm6PQCf5R0
19LvJepk6jsAW8Oe6WQQmeWhf+2mbne9yEsQ7l3DAd04qxfAZuvZoAZwyUDwa+Vz
r7Ap/viBInqWbCbS8W9WtT9X1QqGM7Cz+AkuBnx34B6y5Z7NnfLIO7+ecCz71ZcK
jp51lYMzbd8KAAD7EJ2PmcSLoBsJA8EwELOh90ozLszWfunzWqnyE+govsTk4YWE
djBSjAKdgsN9PdNwwrSTskSRcp/1XmOGD+ja0vV4m9PXGPJpVyiF+f4gdxNSP1cs
TlA04y7CageA3N71I7GSoPl7/7CKszGzWsLraa1jKdB6uZ5sxRnwf8bXAu/c33HI
9vbxbjtm4Rin25PopJPu5njLWZ7iNZPohIrvDTE7sZt4twhUElzwFwCsdztB+aZV
4IT0FqaZF84H5EHxpfQU+VXGfmA6QLwpProktoWq5qe6PRz3G6nSnHCFMkJT/6Wq
QuYrLIluHAjbj1CyQES8W8q2cby3j5iyWjl1A1QD0V5weRm2bu9KJSpu1LXf1/BH
tbGgz7MIduVLsWiPXd2lg1PEqjUQb8wXQWirYnUNYkYcUzfG3M8XeWYA49JbgXlC
e9kNtfnHYmAd7/pWNXn1LD9mt7MEs/j5YciYTMsOKy3PiXnTdiaLxfjCyZr47Zg9
Jg+VBsejVV+J15SNA8ckVVm3qS0JCtyeX0Ey7MBy1EpgX57/q/pUvBa20OE/1XXk
QNaK35knchs+2x+UWB0N5nT8OSaQt6BAE6AEhSN8DUkrrpEAGY+JruQBULsXY5Ha
BcGyHEv2Q2b7AWKwMvz1HuVS6fJymsojtiFg+diLD8ph82if7Ibie4xkyFWkCXwo
WYERsZLHBgyrXB2HdwRukXlCyuM0lBuyFVnDbr/XirT0xxeUBxoRIda11mfOjNKL
+6p0RUVcuLHsZf8KpmhgEjuc/GNLkCyKX53P4/ECjKl0ZMGiC5+Y2QjTUu8eK/8W
hZgNhQoaiIBh9dWrtqyABFI5sW6hVsKZN0sV53E7BGIlyhqfuIQ4TWmgFDjqUExg
eqcuht6sYxvsfJek1Rf27v0K84mu+NmqWdtwCZh5QvrKzCPCijNcE9Lk/e+zW4EV
swnvEAhS5sY7T8skzy+d8BMcgRqZ6g0H5l8FC7vgR30PFGljeSRtm7CIjh4gmays
EsOyoljtgtYOrdPRkl9AAxJm+9lI+3TufKH6cduBrdwl0PknXE1L1qq+bhelcm++
NyuIbafD52L7AtrNZnZFbS7TVJsL7H9VVkPu9yYD2tsK/RxMe9TYcVCx4cMYQFyI
z+ZFpQYxBop8IU2yAR4+f9ap1AkbeEiV9wCJ1FcH+HeJ46mPh5pSqAc9vgzOXVj+
wAyi01ghfRoZqXIZljtDdD5zXAHuZ+kBSausHKuBqzmXTCkpjB7DTzdlAglal5kz
jZQ1QvBo84vvaR+epKKN8EpOMVgAyDS49JE1s4xQVsChF1T9yc4MdzGrZ3EkcIOG
/bdCK9v2JaKsud5ORsRGjwqB+vHxoiWhYxFBnU1InlcVr3TtHcZ2j6Lg4Hr38Y/R
0PNF6N0Hjb3fGCbaF67x16HWCHYujfnYXeSx3DgOaFfsWXZsgfeIywh+vZTzX01z
DRRNIYordkh5zgI9fQ+AQPVf+AvgEy2qR+RJZUwRHYyaOpAABDefmSaKKLiGg0BZ
lRF1IRwslQl+HVVLt93gv7tz1zARb6NpUW+/Mm6sqgkfOCDWsKJVYJHd1EOt5yCG
/TxhavZ5c8VmaEHJ6bJK8H17eJJv5ndcnnni9TTvhy3OQjpyI3EACgeYAU/vZOS7
rX8yHIFpMIdN6cSh3c2vVzGJiquFB5Scj/Xrk60iefUqkGI/HF817XrEp2ijb6xP
eoBzAqZyJ6esypMk37H9xQVT0wWf5gOCaevqMiIcbJ8wwvuOyh5UeNAzuMEfdHQ9
sfObmRDBfrkRj+DKy8qd1JKB5rlzd3N36/JiDYDTI7P4K3dp1DrKQXOcY6N+w/2J
tXikwyFqWvKwy91KS34/bvDEveTt7uPCq8Fs2JO7QCi3qyQuasOQo9U2a2ZjnRq/
LyVhEYCAgRiSCsJDlrcO7OuRu/10r7yza/2w10yeg2hNAUv346/qzO0huaQe3/uB
zyjR+XMBQTjkgJXmw2IdiDw9Uk2sXf+Cd4uvp7eHGOqXfwY5UEox8VuRKNqqhAjA
jDZNF59cD4n5/0xE9Xp+T25b0umm5IQspPdDo5aAKBDAWVsfsgko9qF4dfBZI2dV
3KluuanSR6zhtXyXt3O3aHV4GDOLYLezEPFZJ+lnGFFxRWInMawAQUOEy92lYJmj
eQmdt+pcLOiklnvqK3LBPGuMl9Sqk10R60bw1vBdRT6glmAo+LdDozKvyWzWpyv/
uJSfY94Ul2gyiZPQ2R8l9l0gm8acL+oRIfuQULCOrXVjqwBltKk8+jJ7ML+12RLH
0qnnjz84SY0Nhv0HcjDTgWkb9grxXYVFVImsI9/PFLVrUHJMkK7O3joS4KNi3TGd
KKySzRaDo+KfNEt3yl/KFcWwyAtIlvXG8kvVr1OknfS9ts7IcQ9AW94GLjPAsWO4
+Aw3Q1tk8fbgXILxAKqBrTEWC62uopRL0CCddTlErh8bNlp782KS09KvDAKIExyX
Lo0OAePgjpyKGaoQj50GJEMzXtXoCgUR/HM43FSmIcYlCSYO4Gba7bnEtCub3VBq
6UYv2g7oWp63txutz5dbY156JeLlu3/m6PeG6YllNgqCT3faQIOMEP41Lvbxs7rx
SDJrkewmuvg7VLh9rxuTt+N5Fqc/kGR58KGvHUWa8AqM3RJD8MQRvSVTZqFhpVjR
Htl41Zc6s2eSnXscxuAeMNSVKOxoxQ/kNqhT590RgSBPobo3lyjd71ppzQ+1K5hU
5ya9ZYETfLhgy0p8NURgD4KZNwuDMXoKQJU8yaZUfOFt8azpqSLh9n97uL2G9BWP
7TiYm3nd2I2WNc3zA4EWxoSjhelg6TZpySSNjmaBpp/UZLELS8+XjX8bNAlCcoVM
A3Pbmul0nWbXgJJDGlGzGCRo/e+8AVKFUD74VLGEyMCWUMu5oqmGLldVWFCMBY71
+4p/Ke/m1JMj7+wL4HS1hwTazxmkPki2sfAAw5ZDmNPJO9YwRjQ3Sf7eqd+9S9KS
DFgpTsadi42JyXn2l/tN+0T1YwyqmqfyLXdQUC9Ir2tZAEtsK01nVndeZPiEsKHA
HxrpZpHFpmqUNEBqdqwVp8lk0pEiY1PY+118JChg9B4n8GNLxC3M5oU/6BQy6Fva
tTBDrlsY0ZWw3gki8N1OzmXPFqvOFufVXmhGC10511wnQ2YTpca495Urs5KBuRZb
EMnIII0VMYBbpbcyyFY5pHqVg0IulNYKhVFhptJT0igDPpZPhxVtbOcdOQ1QeOaE
mBx9OJBKMO9w6b3c8NAkOn/AM93Lc7KEHsgyX7tq+l0V8jrby7LTdRjA/GFHd29A
T7Y6VRoWLu7tzzEoqwymcFgFt0mvq4b2JWYDZU1VUry1NT/sKjnVWBebSMeLCZOE
wZ1vaJSDSVbxZpHHT6NZGzqHmnvV73iA4XTN8jvlyuylyUFKNIfJFID56ru0JCTd
J2hNFz0zeQ/4tio1LLXOX7maRMVHItvyrlhWryo/CTm7JjqWo6wy44lxy76DsH4t
HdHgxDUWGUY/1Q+tqjWmKBxD6frvB0nRnTuzgeX9Ll0Dcv2xFYIAydEYiISi2V9a
esOnGk8VJ4Swfzk9ztP6awwzyBWPx/Oi4h+zXQAIZRH6K/uwyXQAOwmKOy5JX6Aw
fw178JjYJhtjh7bU3xzfocqHNuH/opSgtdSXULjg6uTsqu0ukG6KVXvPMdtVHta7
PkrqHar0PcGjvf1qvvWeLSKC7AroIxtTZMOoBKo8K0CqcHfbQb4oRv2Aq0ywxKRq
f/gEohm5uKYCbZAoMIeYHJlBRrroCwtKc4Fzf2chY3oE8EvOu+zhe9BWzy3/ULzw
W5KhLEts2ztmqnSmUfPIeCyoRVN9syLm0alQxVK35ZJEHbBC6JpJBFLsBCY3DWNd
HHSx2KAIDM8xjNjprg015YJ/crUADHGXYCXTyCcvJxOrd/MolKuSXS8Fwhk0VntY
NF2trhx22uMOJtAitrjK6ybe+FPq0bMChR+DQUMtdJVidUA1jvY1jrjriPnTww4G
IHSF/bNb7wMUjOK6ili8UFwb6KWaoMWQadxjZGtKYHY0MRJgQE3dVzOwsHRH51ga
QDpQxgMUcaUGV4wlpP1D/FH6o8QHTMKFDk0XpGPedWG4uevc4Md5U9j1LRn8jjSv
ytm9dlj5LrdurytQAxvC+rDYEQKasu6lnSQtaIv4DDc+HrObYc1IvN0yIEm0udCH
IzQGaFHQgRdoqrkx3dkuTBPVTmp52HkqyXn4XmWQhHN2hX4FEZj+YCn15lETN5xW
Xm25kvIOB7bWGf/JVP8bFg7ISUMmKTRLiDz3qzYKVts2J3YlDpmIXSUruylM13n8
QqZ8n5RAaYn2Dk6F/7X9MUnINR8EjrfuZKqr0a/NjoIrhO8qr/j/E4A/gZsg4d5x
oNGq3JXv/XPwsVz1TAAinP3jDD6JustMqGfXmhTZLixBRKBWXgF5vBgPVg5YuFhb
TWeinnA/Anhqb0ofpDpmqYPQKphBWzXsGVG+X35Jzg8Ocp1HC4LiO3DCma2io0e1
O9PMIy//M4ScovJXYGUrfo52ZJ3vkHUogIdi64mPKzLw7E0jR/cOHzd9nFospRr1
YleDYIhJVwdGMB+dhplQsHvFMo/mFII7wTIB8jHTinWwoJDOgeLj9bysOnmqUMHs
2n0DbB7RqC9sFycXM8i0A3arJIBPVVi2dk1h3xNIjWJOpNOdrBMcrPoKGpdTZfwN
REEVgX8eaP3+KJj7GwyTzItHT3H5OTo1ZdtRUN2kim9MbjVg+NUxQJpmXxhZU0B3
gLyuwHg0ZtKzH9j0DvtmS6BD8WZx+ju0f+tyJ1OrsxCpeI26I2SbCjqiHZ7GuJSU
O3xCHqkHsrBoE7GCRw0ev4klgo5hRHH9sBk/0YsYFj7x1Ie6n96vYzVoKTMnRxQq
y2QgOCVOPo3iaPuUkHzgQGjrhELE1YU/iVM7U5tG636hVm7J+atf+jds5P/ZtTLR
3pzSR92pw77yHY4FYPGyihEZLn0LBZjPOfyWO3S3R/PZ0KrEI0hTueFoCNJSrt6Q
xTzFu4Vc+5hJTAewK+aIc33U1hkjp3kR/ZGXr8D3catGFa3nLfihAo0z4lEBzdsz
NVu/CXOc6jQ6JRADQGQDpTzfseRfqJj0SAKPboFf5DYMaNYvURy9XugDBnQjF2Gf
oCnqYnrE14fHkCqJbpQm2Ti2/1fC2DFg+8qde+96eAQ/GB0/PdL5V+PobzlN1uRe
XfkDSz8I34JqK+TSv40euaAACp79qp+jtj1o5a1dpGmWkDPny6sa0g7MJpKeF9WY
Y6smTz3aRp2o8PMqalzx17yI7IGS/pzusseQlyRDPgZPqq3R9QL0df8hW3pUPNOL
xuhEVzwkNZ9bUl/F/Wvzmskas1q2jXA+ZRCvQ8oNTaLZmLQK9stujkdz7dosMkMN
+VZbLwCvdFbpE56XJ25Q1SQpzkTepBXRq5KVOb4hrIyb+dN1BEy1pXCF8qyfNXmt
2yLfyqTnjmwCkh4AapExSv3dTYo4pCeORCZR0OSNRolTh5uSVrMI/TdYDcy/r1It
BW5IIC8qUYDqu//Ush+f3yDb/lJqQh2fEyjkHC9bhhIsTNcwWh1CTiXjJQcI8mzb
rY6uJ5+97D3UTegfAo1/HWnfimepYEtvqM+mnb6VzUXadaQChccGCXXw03cR+pUa
0UQyAvnUicCjMXoAwEKRi/lN5XsIBE48PiWG8re+FlkEDkr00l827/LBnHCOI8w+
mzxG0HNGWQejZhws14+4x/Y/DYzv1BNcMDQQAUD8aDiwz3Rl5rXWyOiZA/twF1Tf
N0jBcytJi4WiAvAx1Uu80vMQJgB3wU1m1kRHjyoGjv7J/2BvIzsgT/NBJd5bUnjr
Fv4S6uHTpkuedHxXq1Gkb3N3SHhjl/umxF5LmgyvONR9sNMYuA/3KPtnljdlCi6t
2UDSIYufp9vrZdCNxIB5Jg+ts/zyfeS+0IvCrxjYbhYZrboV7X657retDSk37mLh
xE/xl29lteZkRB5c0BlRMbvfReAzlrLU+UNvJYbtXUkzpRE+cbHmIu7F9UecHn+9
JwpgK82MQEUu3FwpmE6IbYYjcZ3OVf2ikPQb47mlKasMdYmgQlW6Cl0QDVNAlI/V
H9S70rngKyyEsFQm7H4PHTgziTTCh/SOTzu0yfPVdLAzXJXCy/xP617XymZBT2/r
ayOKUrrtqsLk9xqOKUPked8mX6NT63oRNgZoOfVraWFIK50gffoEiJD8vsoIjwzX
wskWj62EgJe5sWHfYyTapQn4BRpmOtDmcZX9hOoKLqDDp6n2Qi07tiF1N0bmwIix
6xS93kF18th/reztBy9BIQqfkP9VxQXcGt9qLWwYeogEOq2wjjvC4JHhiIjBThu0
zU5Lco5tZtRCgX/5T8bD+/DFCuRn1V3rp+/kY+qO7Y67PzCJavEx071MTojwtxTe
Jkgo8xtr05FO+3huw3okwuur3q/AB51THUL9PW00QG6g1u4qgoQtrzzFzmopCprK
cMiTThoFtcPauLVNM+Daflkc1Jn3TCKpGU0vpJy05rIORLFCzyyBWJptcbAerGi9
wxd+4QYhUidSTSu+3TJQ3KkXHyGJ6zkGmo2e/0X1PBMNqevguezAP1lL65OGM1du
c2QUsSYStviPCyqHuOAY9Yp3ChNXck1DQ3r2jWMak+YDjNGXIutkPc4b4M9r1RNs
oqDdyIcDTcRQg55d+h6NignjU6na0s28HWjRwHYqbU/yr2lKohnuKvso/rjFG8HR
OeQ0IlyV9dHsw+exua55E+p7ikt/rvV9M3L/WucUfqryVjxd3GcnmvsMBr7zJQXz
gVarvkU/qqubSwGBMtctTcb3z6zKRecEECEg99MfWVwaOb1w4CPlCtIiOFMz5ixF
jth4lHVtvFqWaH0uFQoksiPo8OnT1u2AhqBVal/+M1HSLUCyKVAa1YzSf9xlCh3m
78+/dEspOchAMuKYzzjd//JYaMMKpYaV9IMpFHzo4ZEFPPT9pVeG80VfsRYL/Y6p
u+z6fO3ssVt4j89UKVGIh8M1jhZ6pExjaYCNx0dmE7kw5kBXO+T4vMDl3BZy5y+Q
DR9pCKZ48G7EkDa85CeaX+f+gZ3cxiWR44OOEYtWSd56D/4aFRvqvnLrXMo4iHYb
aU3J2GMsNEQMlkauOBk56ubUryMYDhvzGBzqo+GKgUu7CrJgKqq9UZ6cG9EeS83l
uanqy014ELhduJo7cEBIE76YGzLWJv1WekwEL8NB94zv6HcRVmGB+MmXWVHt2Go7
xRu0vKEZ9p1ajZHqnHlUCQ3tGXDBqrYtk3MxXxLTbpauHD96RkHMzJlQeGP/PaDW
yzXzeYqF0ppnCqdMij5ah9O0cI3XSTeTcORWyGtWPnb4M9Ke5x+uP7UayPM8USS7
7/OtyRaJo4mL0ddUsVNe4sH0iIWpt5RtLkNPc0vMa92LRAHKKBLWUnQTnKeewDug
eIdpg39THLM+cP0/3pNi6uS7mAsI/ZCe9Nn2R+FvvXFAlwxAbxc79jqVUep3wSAW
5OxhYYQNaylCaxLz85E389euuxoLjKCM/+u59XYSZhVFlYIqHCIQkoqqQgOpfk0q
rXvEbvTIisD2iWFgC0bNBhsdXgythXrWOYqJ///gjqVL00XMRaw3SM2AEgmmKhHY
eotDCNt3DBQvCICQ0H5DjyFYO+onvRABQnFCYnFPI+aOoQE1/0lGUzrsxfuOq6BI
vXowoft6GisxPdPEPu1qad6+uydtl5zNMz3W+0MqrXMUBuU4v9bUl9ZKP99KmssV
NZ0GIp0zWfv4BRBARgMbJhrkjisL6xAJniJxFh4qNOinIRTTNF7B7DOkvgnfZ6nk
fP61tg9PI5Cq/zegAMWsH5IawktcdOpM0Vzr0lbCS8R6A9Uh/Frz8j3anO/FHU+g
uWhWi76XftFIBOiGDR6Hbv0gMnLYQGFbdmf56mSc+LE=
`pragma protect end_protected

`endif // `ifndef _VSL_SBE_SV_


