//----------------------------------------------------------------------
/**
 * @file vf_axi_fc.sv
 * @brief Defines VF AXI functional coverage class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_FC_SV_
`define _VF_AXI_FC_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
nF4Vp5YvbO8SRU0M+YYvqg09o+g63RH2EKbLQiTfxqGR1WeTn1nmpDz9TuXU+U7p
v4JqO2qJ8HLe6Tk2ZdA8+heE6lYfTNgF6VmD3cfqSXk30n/oZg9yGpN41GkiYt8C
uXFoWCzsRY1eXWFllneGAYDjfM7yKS9p2qTHeCCrjhUdE1EdVfwQqH781HNhtHaK
jy2D2luTFfoNNAmFQiVGixpO04CAy7WdCDVah3HT8tbIr6HilcNyh+8JTporYNM3
CnHvWjPzuoX56GpqwT4pmNRRvg77t4NK2UkyCkAUCKxqK3eLvrwVatX7ZFBVK3iW
LrNYhykuvPAofCWNE0HITg==
`pragma protect data_block
keu0nc7eIA9GzoSiLn/5SGv9jdLoV1gyfI3OaFxKvJ41FvdIFxrvbyjzktphjczR
gX9K5aiAtG073oCXV5F1OyRT1wb9LYAlnAEYYkiF4epH4JiZuBPUFzS4s4FjteLG
AYbLzkoj1F7+rG7jh5QMuXoAH4J5VdN8hba8eba6W2ZeSsXs0UcgU+gKm7r6DDQL
/OMGN+qRqedId/+tSW8KU5dDUvVRw69F/nIx0qwj7pwBwNb6vxS3pfsbRp1BEQMk
ipWl0m8J7pYTcrOIkVOdSBh0WrYOq9rjLfE1nRCAByrrWGzXb1MuPruASXn4NFIF
y3sj7mrT2dtkspPHZXeaNtZD/xVjnOZnXnCrHeu/HXrpFz9JHOqFHzT6X05gytDh
9TDLr6tHzNZwIb0zis0FzMWb1HCQFHtGe741CcJZvpz4yjeEn6OsYjXqwMLCZgwl
+cGXBkCYTvG4J3hdqrNfxeLYd5qUgjcHVA1P+lyPlsu6W882bYp0pAJYm1Oo8xCt
5Y5gCwkHqa9ZGJpjYycAQ0w+N7wb5WAvIzn02RORYU6jhlo6lOk74GklL3W0sj7G
sJ4G2gKQGIv3H28YnG4o5s5OsDT7yTTxAkOE6IhtfKpNefE0CurHaFRSQMFQDLI6
cnp0NtaUocDyKOpggB2Pv2lx0QTx8QIunwOEKTioD/iX4xSrbfnqTCPiJxlGZNgd
PWFJ7OxuxNTBcB1Nsj2QX8hURW4ov5CWJCePIhsc+2UxudvKXYOg3n/eTi7Or/ZR
9L0Qm9Ean/7NoZ1qSaF5OknJ9OcgF7jgNjN66JVO4fo0co7lzjSo2mprO1c0cLme
kA3vUMUYHgOKyQcGQ83BU7pYTFO/qrtEkfI1A4BjzDH1kAq5Jney2Vl/xOW/Bx2p
pTm5DrXMWnUVhWpA9Cu2fwosOH4+nzm20aBQdgcrozJ7yD5J3o/uW7Tx0Thi0Nv2
FyqfoklZROSSDq9hN5nYun+qBfdC2qhqRz3fWSJQdPRiuzMbsqVwBraYPc5gtZMq
vm49UO7T66/8oCcpwnuNOrmLdlygxBpbeVV+8Vl24lrxaEmYBlK3TLti+tV9KUfv
Ad2wDKtkqvRaEYpw1VGr5g1p2eBy4qmxg+WHUqIZDrNedrGHObgAIAq6dG9AlHw+
TCeMasDqB1lK1/TgNNpNZPEuMesnQopye4lW74QZzQhhCoAwafqQH6VtaCfynoqw
gCICqaW8zYlVlIDNtQriH2XQ1jFTweEHipWdjNXt5LZvJDvMwoxtWhnlHuO+Lyrd
irf6zbdxPRPl6ZDM8CorR1lR7JlmKMNq2FQ9MA/oiXXP6kdIZOwf8Vdlx4xGpFOy
g7vZQhmrI/rr5iLLVlaZmUDSxURYZbczT0RkqRBcSgQy+U+5zlg45jpsYeQNuoRI
1in6lzfJba0GbPJuNWQZUVArQJGnefLWSQp4ZZdHHqnIO95yF216lu9I5YvMwFFV
3/4bB7dTkdliAS17rDYzP1MuF1Jjvf+IzRgSQ3ZaEi5Q8cFWivob3zhrTUcmxmmB
CL39tfQIyTXe36dEHlV9Z2fSAyObfAyOAIq6Qi4BV+5XX7mNdp420fHtYiVQrYo8
D7M/RWS36Fji9eSb+uNUuuSko0+zYdYUd2/T/vtZw16NiC4E+Bg4lgPg0mWnquHR
cey1A6IUcnaZPGrQ6vgt1zBdF4ZBT8E47kEkzm6aGDMFo4CVu6k1GRiAbphSR2Yz
wmo308LCq9ILPAPwtroo+QJiqbXjyOmtvapQpuTI0mzGj8ACPmph0071ewAGEnKN
8Rg7dwIYSGSgWKj+YcWkclO7HeifHv1xm7wTZu9lW2v/fnXOydpTwaVm7droqKrb
6Qztbb4pJKxqn2BUvaMWUX9f1jWkFZMzk2kod3nGouW+eA9lvmWRT/2rkBv/VGzw
NSoQ1LHEOQvokgzf6PzHzozsew17UxuIAiAnb8eDAMczGDDZ+9fA8XgO1+usetn9
FISJRiALnTBo5ynUjGFpKyXDnLt4PZuzuPKsYPIp/CiZnGAq2/PyRUghAatdkbtU
3l7PL3evkeMIczdCoswLqxQCEVIDhBzi3YX3eX3+f7CQ2XXZwoAw6NBz/vYfN35g
WRSecwc0UIGTFA7b3zX98b+XkmNBMADG0aZXEGmlaheQFg5fAyUTx3N0z9poyX3K
bgwJ2GL8JOu6Z7jlRyJabcj17hTIJAUdU5QY/2qHWLiYPzXURLuU39na/TPVsdko
05PzL9HRZI/uUCjHf3KTOEe30s4JIn0a4ZTrnHRXkl/PdsX/Zi5u7UUZOc/5XToA
ORPEFB0897KbIyOTmLoShh5vLs24jvzHLJTKT3FRIe+q7dIwB+YzGv1n6Unp8d8G
u0/6QHTA4cOgbOLBO6Y2YM/NOnVsjgzr6i10pAHgGT2nDMApydOMn4YJ/M4CgDlz
ed37bN37/e8ElFjZYGZxv8NIU2K4u3Wgokjm+FQZPP01ALwFPPWPxpjr8VhlaUq4
R+drFjjgL7UKVAhL9ymXQo3euttDCM3wlF8tuJCO2ItjCDGKGDXLYhAWlrrQH+61
Uc2aRihoZSPMmjwuY/aoC8dJwIKdbV3BxQv44Gzj7sMsac1pfuaAFidgGS0ViYSw
LKUV7eykHeXCNrlkx1PaQ8G/esCnfqge1siN9lkaP77dE+sqUETOJBd3NopowDgY
P2z49wCHMYcfLZIp98Z30oY/AYYr68OJFAw2FgnU+vCrtD6SJlL8+ewORUHot/2j
kF/6bm1JFzjDjqjWQO9zZCq0GZuKFFIrAr3js8IUbMXH6EfmYXaB+Z/3QWESIMeo
v7McTthu+SAYNtFvpUpzKI9x47weL8fstPQEzl2mgezCeZjg5uToDJ+O1jmWTm66
F8b2QhwBkciA1RoLjFbg3vfbHr9qa2TqWpoyO9+ZGlcNfo8DNaHxvo5dTo7It588
jGZNydys7wlLuKsAobsOignAi2OUeIsDNpHuqzOPlJkg79x+NXpf1096PqX03NV5
sUlliAYJ9Yb1NbeN2dmHTuJ2WfroqjkN5GDEc8QIj4SbuB1mJ+trfL2EhBHZqYW/
gvJfSuTiy5DRGrHWBEkVZs5l+FIrAGHoY+qVqQRiFhipBuuUgVa+uVzgCQ4JMHA0
YCylUCuN3uEIXRh/Vmug3L0VPi6I8mRNly8Lygt6S/7TtbJeCuyxKA0hveN5y30q
NpI0ipTH4pRA86yGZRoDsI3Pi66IFIt8+vOitbmDHHSmL25NiJFeAsOUfgQbPhv2
Uio8EAh1BmNFiSdJstveZSCjlbeS9r0EYOw+xnGoknxfcAe/SfrBJp5ICfTctxfm
q/rK6akgOi3l9/8nUTMlcbk/C+4BJM59uLKHZv9/FX9JGz3I6CGheQKnmmatVrcc
CqFrAW2FQQsqGMou7wuol8+9TZKtReZqJdXTQ9mgqx/7a3h/LhqAEnc8QgRABshU
Sy5BJsIzh5WYJBbwDpImRqG8uCjSJ5CefMu9CZDAftsLAsP/069gVhBj8HilO+tN
/AMk9HSZvhqiQc11o7RhMVq10ttg2ZP9pTFrNAnO4ha4TbLtLGDjUFhTMsiefb3r
D7xazZfolwkEHq3fSCIzFCKw7mLENp1Q3ezWSsa1v3zMr7Z7Lj6ZVlMz8p5GOusR
qhtFjrnlTQjKTCAVyDRiiSi36lgfgCtrOgB4p+bGNjidz5SWXLpSlUu8rWamnbmk
iyjUL1Ea97lkOOttIO0WW1tqi45CdtWM+fu/rDgp+HLiOq88hKBeiHPbVn/nd1Tm
W9TbDpRv1rl8pEX1mdAU4jEtiFnIsSIlXv0s8bwVucL03qv9SI6BDQpoODr+RPL7
5enOaBoll0isrrI6IveCz0Hjy+nFq9ffmXQUm2BnXe7Z9Cyx2t6twAEBIvk9HIEr
4WWT3wZ4F0/O8XOe0XP34A3FFVe8TZjRcUEzsZq/4UQVuqineMvaYcEWxSpHfNbm
jom8mLE9Ivt7zkjlxN9dBBYN+r7MtrHjwUpyPaiLk8dPjjR27wJFEdQxeWxsGesh
IbpSu4xIIPjw4FNvZmTxuwDeqi3eww3XZzST3G7IuVm4QnEgBs5IpgubzhpEN0Xx
OWQwZUvQkhFQ8UDKUUdzlwvb+0pQKij+7A39P+laB78CzpMgihsh7D1D5RFOnc/Y
ZxB48r+P+pu/OA67JQNIEpcQzDrfNNXSXpIbQmjngwUJqV276m+zf2wkYLYstR4u
rGd5qOJq6MIeCvKLxTgOip2dycpq6ioN2Xi3qEkZpqRNieHECP+yI5JsIMfwNnYr
mFaIPv0qHcbrPJvEU2j/RDXSymdsMCfOSyoQ6qSZkwtFV3eRjsHfi3Nj2LDE+OCW
59N2T/4XdBo5fPr5nye3ZhLx/euNlSwXxG96lHHxlXOyO+EUdjkBXyY1RDXBnc5g
WI1e/aWrcbgCb3tdtaZOrT527I7uNzk9esU+uALPp5erhx/+ubS2vw7pV/ABlSbH
bg+zQzinR0jd7TGIXhX3DferhNf9b+alIEXBRm6FpKWuSNnW0meAcf7b5sX8xpc0
J5NwM4Evy42ljRY+WIPIRzb+1IjEVidEjIM3wMI78W1Uf3gKE6griWsAtt/k6bH3
T16Ve2z0ruAV6kk6ncxEFVTgB6eneoTpjQKozbu9hlP0xxGhEe+jN82FR4WpPtZW
+KBBGMzvoysOJlmxJ4IwvaE+DrL2glI9a8i/QfG4Vij6zj9lSdR/uhF9AmPVaJhx
+FybCdac0KAV0iJ9OXvD20JzFvy3iQItitxVgyApDWvCCK8hmU9En14FjHxwcNaz
22ZAD8JIE+/0fgL5sg2pYKTNh3d67D95dNpho6fsor35rbtwVhtnecN4etLeR06U
o/jRZlsZaiODEANeoW4Dvcq0Jhb4Ii6I1Xnh5LzXpHEELQ/H7LzbyYABHoKXeRf+
DTsSqaZwTBhJHQlI6nC4wU1Rel8rIsXj5egBknuT1a5doAKKOjtBju3V5zCSvCVD
qdxevGUjgPZQAX/iJcSTaliAo7zeLGTqkcAnDT95y2Ngk1FpFdffUHekOJn//2T+
47HvyGE6XZdlY68qE2Y7B8J375yjCfBCLRsLlNcYQBfafKy/coH11RBhHseyRSuS
kKkPg+fKwjhh8fQpIahBrovYBCuwxsGcC5JXrlDWzHeOdgD2OAKP7wKE109BjtXv
nL0re9qtz5wZ1ZllJyU/a7EIds4rCFt+CqfIjmJlEYYEnmU6jyvdrag7KTEaImaU
jDFjQLIgsSut4NILaLmMeioNH7zOTDtXIVMx6EGDQNogALtdn9PGEs8/XG41sd2O
0nkzc6XgL0dQRCEW0Zm824hrXuav/pVBQpuiDZ1Z3QWhojsivwdJAvBguAwVrnMz
ARsn04LAzlU6pJ68lAvPkWKNX0ECjQmRan6u8IuiOg7yHIpziEuTvPcwo2FTrT3l
s2CIukwNo/n+JwAyJrf0pdTv5RM82MxhzStc7UhJ4NDJd4QyKa347p1EMnQdrKH/
R4v5+CnAP8OfUNTcqViLvnorQvv7e/+7FswbImx02hcYcK3M/gFPaqhw2sMOoqCf
eUsnaaSJZ9Ii+yLegTzIYga1mPSl/8I/NSS/PiKl6iWQv/mZVgnIEZqID59n6QqV
DovhET+XJ/HvE+g5t/eL1xk9rPvCo2nryNGOj7WnA7eA/Omp/wvrb05wQKWasAPs
Hd9t6KR5x9qIn4Rn0LrRKaxudr2t/ZKEYXbpAnYSdiOLQNTsve1J7frikjFMazp2
d1qlbuIuHUfNPn4T58yqU/SeWS37eN9Y/vxoXwBI/jadNT4gYmZCy2He90SbsCku
2LXCs4jmhuBhjeu7dizT5DJ1elT/Fl1gXukRefE05bLRAcdNABXn5fnXnrN7xnNJ
e4eeBKHHJyqLZrQfAXzdIMEHXRUB2oPufiBNjFvtSpOdLCpbtP+HRvVZutGNLP+4
nJMYLEAEWlkqkPlgJ9AP7ywSyCSWu2AXrWPlCcigzL8y6fUr+JXOoVVaHecv4N+y
CnUGc2y0/OneDnjFRh+oX604egSE0R80QEaioOJC/ZSLyixh+T8A8l8ekSJ7S/KM
NQlqoGjNfpbbUhGgOmKyi8cZji43FAwohRf/5opuNQhrgNBuVqheJVHWw9ZlvzNr
fU09hG37RPndyX6fe8NF5TXxf/mfbpDxekR6rMUexx/AFRQzpLRMre68tkdKqkLa
gYu2x3+8rvB8F9TVoqwxzL21rwqZ1mGs0jRhO8njjqJZH1rfaKyDKOxdlOn/7e4n
Cgn4MNWE4p9dsJojJwfDOuC6ZZgHpW4sVgiiNLrlyysobt3nCUDwPWPPGxlxwQqS
0nC9/4ggwZwFo4eKHj0I/gya9Nnoe7Cz3K+XXz9LaDyycXaBwqulSJI9C3xrrYAb
Df5S2ZWErn8AU3th0egDiVkEuup+J+9pn6CNH+BglGkO958FitEXK4wXFWym3uTE
g4qcUMiORvYgeYbvpcXE2w10w1kgpQaTumbInGdl6o79IiW7dl9R5dBYl15b2qbP
DjEXXGvVXRtgHPFYXs8D7Ojb7+YKJUlf518Xge8HzjepE5CrEM3oeqMzKaASQaCp
5PTZId8NghAqrGH+yGZk0L/GWCireSHe7V/Xr0QcJXu9JMJP5lRK1HcFAx89sPlK
uSjgnkCBPgf0Ds6ZC9s0jJi0pxQnhKn5jsoFeC1rxOiR9VHcFEZ/RwCYzrcjcs6v
KAh6YqA3tnQI9Rk2CTNOjqgmYxrR7mtwi5VoK92NnVmme763BxSFWkslVNVHpkx7
jAoIfvsV51oqNcljiX3imayp4v1W81OzQT2/5R/g6UYfi8c9lrZSJ51vIVMZgolW
HQPNVrEOKhN0157Xwwrt17Hzu7TcVw1MLnK8qy28XYCNGegGJfDbSUwCFVFp2hzK
J3zKKeoT2eG8oYt4uwldXOumMDa2NyxCnQYtJypZJV/CzSnYRmvBPI6be1CByg8z
1Ps3n1OS3e97LpXR7Q6BBdNeMlX0xwM8qiyLwbv8zf3bQJO/GzdkrPCXIkfVJaGr
+jnRDVAtmcsPwgJl1g9jhVyqCC27Myrsd0lx5FzvJ1zwTRwJzXhMlPq2xu5VqT5c
C1DZ6juxtTdMAC0TY5NRa3qtBac4MdZoTH+Ss7xovdCQTWXtwp9yfP0441Q947VY
ordsBaaGFEfjENtSoNjSRyZPlKtIV+mc6zCYSKGkP0KALAwEbEuLluP5OX89CnPa
JY3RRJ+yQ37ir/9mekv3mckHDcRNyeCwz/7O+vI6nvFuSd9UN4vnPfh8H+OnTmVV
+YGAoJ/NxUXS1UEC4rGnpiEsvTyexMAAeA+2dDF1erTO17dT7yFF3kKIUg1qwfN/
9WrGEO2oXqMqkvVyDpU1NR1/aqQmnCOiK6SOpRPEGxOoLeXdskqPVC/XEH9kNBlV
rIBXbrnYtiYhbU4WT7ShzKvqCVjMnIZRH0y2+T3dPZYSgejq9G9Yb/9HFiZySUNc
1djrrbSLyGIUVzPDMI9JJEWPp6v3pj9iyirY9zu/ybmBC1SXrl/pBZK83IKqUN8R
VxlAhzihfdQoBgR02gQKTWPTCqLHei+aVdoxxUCxaPqny92Rm/vOvmDb+co3H8At
vMWdi0UWBxSDGnfwMyiqmiBJBdDZNRcHWhUChsAtn9RhlGJRc8dy6YekNMQaSAhJ
ZPKZtxw0L35scETupxxIyy7MV72rrSCKr9aJXUvNTbHn/6bTkXam+5zKKacSON2I
A3ukOHzcjEeBTbey/fnXrKh2DEC6L4uEHzuxMxh/RmCm+4mXU4M030hUhWvKHQn7
EcIUmTZ+eXE4V21N8OAjweUmKPUhzywwEeDeOpErxEo9CmCGqyJSIvUYVcspZPBX
PEtdPMbJfFwwludURFEYv2zSpxDKOEZKKqGOc+PIeuz8rQ3DD8wAKGcknK/HOgN2
DFjlMIHRq5xDr4CgYMo/u0NFPD2Ze9wPgx7r7Em17t9NqnuXic/Uk7VvCBPU1mex
sb3iGhpYPcUufHtLgD5ipEQ6hyFYhiEJaXEiAiOMJs1Cw4lphzrSsYK0xVpgPhoL
CMcPVhTfR0oqhFuzzlbFkXpYX2/Hlgqa8Kn61YZSNUlP3KsYJGC/vpFSTErm7Qvu
OTOv9GVhpYV9bLMXFv81W5qifZ3jWDrTIdQqwnUapuwpp1mi8uxZHKYgyhAqR24x
ndJWDc6PS9DP/FtxB0ZBUiJAcmE9P4EDllETUYvZcTRRltvAjW1R/6bmLqXQSkGf
sir3gzHlIP4R0L+j9/ZIx04pgbx7SRBkjYuXOHOxzWUQlusbmiMV2KaF5OjMtiQE
CFC4yxl7wiDKAPOIlScJE7EE1MZsSKVM9nnyT0VqjN8XW+x9pCQIEgprPtqGoNRN
4XhgzWwzq9lCizJ/YnJ3Q+btiD0iP9PGpteLboAp8vaE9v0Z5ypi8Kx9kpEV3x28
7DXYcbe9Fqyyst3xBtWYoOfR7WyLUjU0oyEweWgqYaayMviYEOh52J447lD+RN6G
2I6HTvCRkKzxldOGJn/c+kQNvZTn1cGhOOKQHfmIWA3vzf54kWr2bXXUt9Qu56bI
t5YrB3MLbAPQyh8LA6Z5IT6psVykgH9hB6kudn1cEEUzYT6WGhNz/RGWFCS/Xklz
0YoEPKxTvD3MEiKZYUVlXL/eb6Ekk6NVJ4zhOZS5bDTre1lVmlkpTQ2AhnW3Op1G
Iy/1NPtykMUJVzg+FUQIvIK82msVSaKGCjbjIiR0jYCIzlcplVat+qbq5pADiZ3t
6l3C8jocrRCfDK7PKNgGtxivbGgWqclkGEgB8V1OW6VxgZ6pR4Tceo56wlk23u0z
t/OOvxKlNkNqAKlJvBfIE930mmsvebG8aURWnTXuk3iyXlONrOaOpSSD7M/bO/An
Kw6frjK2T8MypeUgcMb3m3oVWRj/oH+NyTTMw29dFU4yx04FWT03HNuM6HCKMPsP
A7dRwPrSadFRSacC/QgCRYHkOAEJ+sfh8b0C9BWftcLPLBG1HiSLeKOum43P0Huh
IOu0y6DZC0TAY44XHaVEyiJGB3kuje2WtlN9cB/Fb9jPgA4X/WngiQs72sLs4R7G
N2zXwJriXn87PK+69YwoJ9rjpUFmJKLqwLKtARNAkiF+tQAWBb7IO0nwE0QUgry/
bgeim5MeaQSsf/Torv0+HNQ2PmYANcVN92TF3+hGEJ1GLnn6KhreDjkZeyzKB79M
lrQPDW4CUkLrAw8goYbHwD0L6yPqkV8RBP5irVjcUYNGnLtfYYbBQdD+S1+ratPj
nn7bIRx66CB1hM371xRmN/sZPdW5eM3IKvkoJfUg6Ipxjx+JsdFjkLUvbyjHyRfa
ULteGStodjbgbZ4L3Kp9opa8A3hdWiPAEjcMau+0SjZc3J9ATuJ1zJCqJWfss/pS
whzhvsFPlyomYIWjcjYZXarqZ5X1ho8NNU/7CsJd72pqg7EVRkZ8FcjoPKyKIK3o
m7Mq/usbQfWr/YtqWJpAfkrzo85tI3V931iBiiAdmGyl1EZxokP6rq5ktUA15txe
hnuM140vgzA4oPHpxzNnOdFyzKlrs6RhvZWZf9DPZWKDUPPdThhh385EG/1DDTSY
LlPaK+AuVXZbo1xf4jitftND5EWD5jNZBq4+tJlnKXoEB0OctLJ/uuXogk87l5PZ
j83iwu82BMVM9KV/rwAha8C8bASLxca4Tp6yBQbHpXLhLoVGTwfPedq71nFeCbnO
2UlknFvW51o6x/YTi7TnrEB0z+397njPfEG/elIowFtpVaHJHDM5+NIC/A2movTF
VBVgk+qP4r1zc6h3Xsq5/ukKCrAmm8tV6tB11NGk1A75AppgDvqkp8TttOsEwXmI
10DNdq3BUVhD5qXbaIW+MsnboHHmAyfYxYgYgKJze9Xq+Qr7qIlVWNazMuq0GBzu
6k6lm/leQwO2t9T6VoYSijqNfq8hfaYXY8aIk+pyoW6NZnfXej4E4Bj5UdGQzByO
qR+9EQ0EjsNEUrNbqTh+5ZAMajIJO0J3Z7pq8tiMbmNhJxE+uksrjhWf/HQ3AN4i
pK0zT7Hme6ga2k8ut33F4DjlBM/Q6JTvHn3GZSwsDz0Y09/mKkBCFob75Jj1sU6g
kcqQLPKj8oYswLQiJHXN5h5iOQ07Ibp/fgn+uiRKvznFENucisgpljEbf88ZYnAK
3n42J1uX0iB2AHnDOo4lRXVxP/OBKnnlHRpWwYnTGKzX7ULTNEwRauweFscy8UX8
+yF/gHv+olEMIZS0X1pce7500xQ2qkfJA/Orwu05HXxVhtgyWkQgbt30oGKGVITt
WnrFbus8Z+wz2gAQ5mufQjnOKhrjxbVLmItABdK+iy1WOwZJB0B3Wg1hTx00/0yd
QpvhZWfFfwMCyS+UqK5FmyqjiExnchlqe3HGWwR3IEhm/bB6EVLKbOH1ElDzxjiU
kfzXhPv0ydG2lvKiI2Ke6bKeQBaG2nT6b/xfONtrPxecByVd/l1NnoKMrJ6N5HXR
y0XKnhov5MWhpFCo6qUfCtA3vF2T6c+5QsWxlw8ecPB1axE0MQL5eIqUEER4wzRE
J8jI1skgDcBBCBHlmmIfjj8nKzu8NDuYqB0GWbanESl4IzYOTC2I4W9ZZ/gSyiXX
2buC9jTdXdIgNWYAhVClmqBwEGSq1JBqwpWfB434VuAhLxo8gZqmRikQ4hSHJhu0
/fPVmI7YsjLlYIPE8LTDq2icm7ZjuqQaRHuu2ecQNPc/IiG1wa5q2pSESpFPJkVT
Tz0naPvLo1VMfWcps3TAvda0wR/G75hTUoeARkhz0zKr1DXyzLdSDOiiKJgvKraq
8ew5GKTqhCXokzHx+vwVbN2tg2LDOW0nFwnF+hOGM3YgTZxv9UlSUTmck9K4Lpn6
+m9h0K80OLfy4ddBNABq620/e8b1suFsUXxMGaTurgRaMAFpQz2l8lBGbsy1/SdL
41eW9a4crFi8EBc2ErYjomNzhnpX3QDHFVbcuhZfblzSSESFhpd+MrrkEMUEU7qM
UkqEV8g9z10o4+O1mcL2MCCZcJa8kspuBP9FHWdauk3B7E12Q61bsfQ1qIGdBBSX
6zg5+rvo/Eck+qUZbs23m11zsDj1O7WIQsLEQlH12pyfA/WWwuBXuAnA4ezD+Z/M
iArOAW+bkEOM4ZuVa0q4H7wxkmBFZgWyOFOPFgVet8SAPb6dH2WkFalwvdYECZPo
0UrTQ0ksfa4b7HINIjDLV+alY8a7oYALBAAjYulsEAc0C3g54LKg9WVFNEBI+Bad
eO4JdfF6+RTeF9p6+XhDbT1Vh2Zexg0i43p1Oegm9ENI7FEdVDjE88HO4911rmK9
jY22G7GYKCLN3xYKxcV/02tiZXIr9I2A41aaGlquu3yA9tYg7KM1UmH3XhsJhAWS
4aUVlPOdIArtpSl1tyJCAKE+GAuIDbjO2ncc+CjRZZx2ChByhLe+GhMGsqLuLzdy
oZqoOYhdMfjxvXHv3TYiHhEuJdv+RwMi+q8V3S9a1T4Kem9AX11la68HCjWaVjjH
BbyTARgQSZMuy1Oy3rqLvtDXkD+tEVTQ6aAUAvLbcxjNyYyT3/m7nqeyM3TMZAxA
m6vB6dJOI/oOeiM3Sy1iVdfSLO7I2GTX+sHtfuQP8uNzrJFuVe+rd8IOOWjOuPGW
YfWaPRB/eOBzp82GnOPySoUJUZs4ObW05gM//txy5dxOwAUZWaMW7dcG5Ep1zrmI
gfH6z21tekybz0fA1DG+w2DKCHGPbiKrF6tb+3DN816qwhvJkNcgqJkuRQTGuAjB
p2Aqo/m1/ZWCBcQO7wIKIA8irzDRg3OZv2qBWYW4BpJjDsfodTZoaIdi2mvk0cee
/G8FwOOGlTkXrlLrl1oEN0yLVhXWqm1eW6a4MF3buLb28mqSh+2BcMG9Icbtp+zt
JISVaRmrOXJdGliZacR2Qn0l/+oxpzZEBgJ1t0LpPaQnh1ovm0nlWEfrqVQduOYI
2nHVz0rCeVsp11JssjhgHScSKcM+8vFrBQjA9cHuI8WIZ8rwupQ+TwcjlyV/jdo1
6oPAYIiPsXfwBrMGEchOa1dZjPGbcQLBmHvrDiUZ3D2nfMeBn/H7Lt6HrZKsxkP5
JZW/s3U32S/m3Jf6Cp/v1nK2DV0rUWWzgphG/xRLk1Uacrld+vPyrwe+c6bjgEmu
HkQ3mYgWGb0T734oHIXvERMclFy1Pl9LLrsb5LzLGChB2Y99BClf4IVPpMjHSUP5
KoxMUI/XoMwcvCvIdKnsiKlNJt6uxsywr66a+vqLFw8sB4torNMKLATtnZfk1PBz
85EFbpypnG0ZywaDv03oiKgiODCYXGpk4Nk7jqMOXe5zwjuyTFZSp88nRJWrxWiS
9RU6vKIW/gsk/D+Q/2gMXma/qjas4yqYF3GoCEF4KmrrtEVFaJtbeCnEQ9n7iciv
CadIX/sLLGN4i4EBXrOkIy8w86yomu4mWrgn/bBMtfb9UfMpzITDsV9EMrpJftSl
0gEFazoCvvUI42Bij8/wwOWnzJpisTA9zAaklnSfvVsb/1HemmExPniL8HS7NA5u
DCW5LFNGYApZ1dIZvaRZ2or4AjIPrzcxrh3bj3plzwTtxhk+vlswPfLjJys5ByMr
4hJ+RFOE06MlQPT9Jcje6/rhNczdzle/pyRYlOgl5gXwwvA4mZTC46hSANEC+4UW
VZ5gPn4YEY/UV2r58+n3MCrVxzNSJW2YeKnNp20fh8pNJUAFaU2fvgUPOAVuJvUz
Nl3FvYQ2mZTTg6x7V7INWCF9uqc5Y7wyniyNVhWm/znDcpLoZAnG8WxsUeETzrkP
bHJ6QtghReuz0Brjo+IOSFxGvmHOnLLAEPNwZ0YAice4Ps7UiF7V7FuSH0DRz/F9
CVQb/iIkuaviz0tjbO2UCwWhfcAyxoe75OxF5YVhWKWzRGGmPa/DqP8hOxNj8uRl
gi1EoKMMakF0kai7wtlD+vFLfUgJlJYmRuGDx+gfgVNgTIhsJmvwIcAOjIP1kRYA
/dEPitwf+lZ9tHF1wHs1VpFqTcvzDMeiI0JNWh6YLjadJshnVjjrwo1xRquZiVQJ
7smX35mWazo/ekgs+Okhqywz6U6m+gVuHKMR709C/k2MPdJPcFeMP1SnkrDR83LT
LB0rmCozr1iTiG3Re4qg9jGT6Hf2oD08fG/sj9Vl3v2XiNTkoM44kzQtXwKhN8rF
4rdOJq8w0K/mHYlyfqCAk9uLZDsCimkevI9NeJwKiqwBvti+8F3SivCrM8qrQZzC
ABnjkRGXjupixbasDoYo/kU4ryMMEfALI3EfNd+gV5lh2yVpOEMkTJiHOwUq68Vw
0SMFOtzZ1wWq2jCvF6I5e6Qthi1U7EJX95evyvK2MVrQ3cwLIlO6y7eCcBI3knim
GAHrfM234l8rCOznfttta8tsq/asbpTO/fVVn01qNUBYxVC0jT++ybjfyTErAwwa
9UHQPgVoEkgfJjv8bUOztbBjvV4zKHxqkcl3yZ9nfvi19dDqCZ07yQwBPrUuIGHW
v65tMR+WCQ8f5XDa0KF6u05mrmHXz8xq0tQpNH30sZQwOk3AjBy0JM0SB9COsH7J
vHr5v1IfZCpLSEEH4Nhngs2FC+iZ0rmJ7dblOtKKLGeWsmx5ZoFJLN7h0BAi4Vvj
TUMU6+8/fTA1cYAkxT342SMJ+RWFzS6L2cQH0NqkIoUdn6bQVBo2ThcosISpn/+6
jhNwcMag60RDHzf2CXjUJ0NE7jUBDSDX5wGZMEA6O8K1svjhj+cO+haF4VbFn7Sq
S4yeaRK31xifjrrNMY524Mfq8m9jVZQ9sk2wtWC9ElitR2QrLkbvbvH1W7NyZjYc
NMDNqTOU1dvf+eDoC30oSFU906zntbAkcSPBdrNDs99frxp/YQjIlMTXVwT5pXiT
v/WC31Tikd6Q7WD+o8zMTBETdj0cBzyxIU/2XNAVtN+ynqixYPgdyP5WzvP/AZBT
9s2xQPdUgNS4Ym0t9Z6RbzXZZFSeBuceGb67NO2/HWliSCxTTjjCPdJA4ei9uJEX
kMrmYCB6HJztfu3+/1p8el9jh7NwyY/FbTq6wPGml7n+ZXJVSTGyJ8RG451AfswI
TrzloD9xq9c15xhO9DtnjlZfKlAk+ByAz1QfFuz5PvIdMcCGAcreFxAiYBOTj7Lj
FXX0eLxF195SmNXlXp+fz6a5i1fzYW378ho22FaQneGZEynJb0WfcWvcCexRA/vA
oJNVZDr1+RZ1ScPk6Toknfoe/reudguaGZqpHthoDEcNKIr1ExWDPXwmOQuSQI0U
4iPu00udmBvDrdZqUPWBLwRrEYjHtqiBmnYIkPEd0euglyOMZ74J210pLNaHjY/D
NzrP/Bq5OLXK5nAJ0jnmXabxQZL8MmCqnEUrggbgWHOgHW8e/XcRDqCQkIDAWJnF
tuMtanPSWQRLX/qo9QDclM9sehKIPmWPffZ/AIgyN8syA7l29nyHfCCO+oCLv3GW
aNTrnQ32pXwbF3vT8fHjl/CfKAN6njqua5AXGNGr8qd6/rY7Gr5zBMV4RlrQ9rYn
ncuDJK8PMIGfXFEVIbP/FzFIPSSyI/QEwUp8YDW1HsRXvy91lP17reecGYdW21w4
Y0XiYPQ9EwTuT02w3UNWb9MBzj7b3ojHsmRSrrxrXtwK8GVLWoeIPLwVfJ3D/QAm
FlbKWnhT/wdY3QPvDwTkgVc3minkObjIcxuz/ICymsIk/2M38N3VRVnsG9o4Vo8N
zxgf+634I22D2DKz1rIDiwLFo2Qoy1+7y1ML1CeSNdiXqm30SbLWJF1bsIF6WOqo
XSc34Ty+DMiDV/xBFkSLJTPoj1p3Z/1bFBZVX68s72aAkQlSEGgluv4gotwE2WOV
UaaBOGv9ybBPArDa3wod69c873XSugIWj6PceID5s8/TOjxXJmUnKF4vzXTl4jfB
PflWKDH8YFWOz2MKlJmzgpbNqFJDTBWLfPuq4ou23zmjyZYW7kiOtSeeu1OyPJyr
3IdmqYetERA0gmYU3KQU3xt6Dkkfb+sW5C+yEVbDF0/Dy4dU5Zv3gb6qJcMeAoSp
d8NpHWAMFRBI8tR8Q/qBn/QpW6pJ1sGF/KZ1yfo7iefKdu0Qv0Ho7rWfnRasz5A6
dOVyxhUnXWyyjsA3iyCJgRnu06SB+4ZfnmI5jljvm9xhR+ErDt5fz/axQygYlGsY
U7myQnCUbjFs6pbCOtidjZ6Ee8J6AEIm0nsMZg0fR0CGhC4b2/gHuWT78IYbRVzm
PU4GgJE9xK92RrfB6BBGrsFF3Rc1p9h/EKLxuGPdRFfa3FdHoDAu3PToeeZn+A9y
vCXi3fMeHANlCMUG7GvyAX8LsrTO+hHokRpEwLPx9Z8VkVvvCmu2iguzhLguLJi7
+IoVCLRQ1mdGmY7ZfPI6qVX7tQMA7A/bQduwurdmZ0GPrXiQi3bndvK/fdBcY+O0
Dys7F+3PzQKMuztNkMGuEavO9ZoND6sBzCtPQg33r8PimoBiBV7eOKOCHFBr1uwz
k5OpWv3QgREh5GO7It5qurvODcYmwlJOSk4pi6jQMipr8O3JUUYt8TjYUGGNm8h8
prwSlEu4k8c3+5XXJVzfvZj5TbxPWGOFVDSAN6DmkaFya/RZl0eQxr3ZyozwwTWy
yrJEyIdgnwKrvmtIx/9ODVNULOxSDIOyjC64cIdn4TRrLWvQ2+Pg7kCD42nVm0HA
ZLo5qU81CpE3ciwDMPlqdgRnvN/I+8UkLlfdnLT8vDLT4YlgoGQDMofAz+AkQTiB
VBDsgkbBkxdWrxUGQsfkfWrsizLQVWwJch/qHWAhJXnVdyG5tHNYqW+fC8OjOaa6
Qr5ODVJkHv10DeQ21akQHWYhbn+jvvo5XP+KTG31DhU9hl18C2zaTdL1Hs3xr8+V
qOgd1Chw+DoYnM9M0U9ghxWe9evPceGNr+gTxYksIsOLfvMSNObXTebwIrkYRW+L
cVEVfbVOL0e5KuOwHPZfNfy3q+hcwFauX3Cbe+/+JW/42PjzUmopapxYq5eggz5P
ZivJC6Y0UIeuzmOKsgdyjs7C85hm68qDG/88FsHyfhzMTTmNTLrB1xRi/zuTj/Kv
5/vgxPhg1z10JK+uU7areX6ZMdoRSIolOVBpyFxAAEWrOWTq4hTEsvkYDuBYoAyO
UVudtA9NMmeuJ32ZWlzTP4gDrt1FFInEh9ZcSnyviXzoZQRVm8XXEMy3LvI5tJow
A4lC+BLRjiQ6WZRbVh5s4evXEB5hz5wFzUjqO1BiRBTh50MOJI7B82eKG883qZQr
ZDsJeY+VMUXCqBlEgcJlzop5LOfYeq0vJfpsS/OCqgzY1WOTLS71sg+jKaKNg5LI
5nII47EHcZtSJQM+AQnJjDaq0RDPSb4Umc3sHVuNXfOcYH69Vtg8vq+G8BA9yAvW
B3mpbw9OB5NwxMwIZIhi8gFN7Q1FSEYZ5ubT3TRXkNsYR2p+HcsbzVqqTXdEl1jr
l75/ZDqy9fe0DeiRk0Gv9ZT4mcR7oU81ciL0O3kZtPlsXQt+k3eBmy/OI5q6Om9Y
qCpnokU+qppSUupQv9fRh2RSJRn99pK6RHKUqcbIkviGwNxOotgPDLuOxnBUzw1z
deVU61j50QBmM3XF//fS/bTnWZh42HHNKDY49qYE82pfoRWXCFZKkaO/0gAjp6E4
L/PQZqIyqoJcgURcKdnP7NFTK/KR4jzo9KtQqfCwKMgEOcb+euvTMBnvt0T0eXCy
6OgrfkvPUsnnvXvmkWzOsaq5fGH09qp0iem+Whwe9IyQ65GRDMoft0tbTFg31klW
B3yJ+LYi3Wxd3MMdxIXgrRz9An+SHdQOciCKfZ0/cObSYx34B7s1ocjWiQqLHq6t
wzf/eZYraoDDQyy2G3U0Vot7XPZiVPOcNYZ6YbEFSQjESDVdgAXEihV0LB0b2b30
WXTExG0g3Tbu5zW24LNS5Q01efrHTeyK3bOPqI1RsXcps0ypA7JvYOgUjoz+f8wO
LjjsLda7pBO2Xvs1nxLPsvDy7vMU2zc8bXujNfl8tIs225cPzogjBKHwkD3a9THO
SGnMRx5e2kb0Y1usHD38uy8w1pRltBfyrLLi1DOZHaFjP5EM0IMe6L/BY7rQ9Siu
WWmrGOBKT1BOj95YTgwwT4Z6C9poKCtlGq+gJcMH+PIK0S6TrHgM9juakqxKDR3B
f+2oqSJuYydLU8iYSmZSR4G1nDfZ1bLJtKoyRikUQi+txqyuH7MsbsTiwt+CSH3e
eZ964IBQhL4YVjoXj5crFC5Pchtj4KgVMHTqtzSmGOTuACLS+Bvm0/Q/f2V/KY8g
1Oh1jCeZrpwsMTTVVEeDSwcvrlWfYa7c2Wmo9zQbua8p8+iHHdt/TRRB5VLlaAe8
48yXZecmS0FvF8dLBGQdnqDr+QztGMvDymf3xaJHcTVuzZZs5cGRSxEkei6/eQcm
WmicTBEShjtwP8AAWai4+rEoyZSU2o74XORs0r4vJPibx+Aplr84hPBfsQEU9R8l
Thh7VvvCrX8g+/34OJVddYRJS4HwZpmFU1eCweKU6RZrkKi/97wka9TKUl+Vg148
PryaiQT8hCKH8DnhNyQoIfoM8C2NkeXHxFblKa9t4DB6y0ulCizLsPNC9gscDmDg
YSmEcDqn15iplhgYRAot/zAKveCXv8LTk4TtDZKsKvGWN902+CD6v+dsXon6OQj1
vSS4KlFMZrMjwzp8tfD7N1HTrtR279iNJpY/vaYPTqDeTMCgCSCUuNcy8DgL125g
PnNU9RN4PCG61GsQn1asWDDUQztdlLoDubm7ahIDslBsRUzEE2R9DHETXWc8eRqH
2O4F9/cJDw3jAVezVHKDEhk/FpeZZIJK6cq9FpE2SDoEeKAvPbjKhO6UJka+eUgH
hWJSLjoM4bhtE5vjRqasORX+68en2Xa8b3D64wpU3hy2ypghdPqVZX2QsZ6ov+ux
wb2sdXlLp9uyEwVaGobTbOWvqUq6ruIPh1F7uTmp78EaNPKDzLQbzI5TxF60/GCg
xH0bEPgd3blkjUnX5kZEVB0gg3M7iUXBM/dLv8lKt5wuTm5/7STgnmKIzvEea2Or
VDbwqhC4VKqPPttTcsrf5172LEHg7BPIa6SvOm5RqB1UHx7PgAeShcfY7bXRqDLN
wKDzDJEoPYlj5ZUDWG/gvLYvZjV9H65idGFUTrJOh360TXV2DL5TsJRvxXNCgSub
wlXvv+xmnp3CbqzTuRKyfOZzeg9b4OtwXbFXlIZ3+730R4zowIY9poZ8VaelMhmk
RJ+nkFRXUMNaKJvcNSdqeARGFpA+PM5Gu4ydiMqL7ZtI4TLe9teNS0ZNzh9bs9HG
V65Asg+eV9WkPZvPR95YXSYGYf7F1sAuzgQVBO6XWPxvosvzRa5vR1cQzmhvXijX
79LQEqt8qSSgsWPDeqxp4tWG3E8tw+w5wBjbiUZI3474rvJy9yCcpcQr8tiE1d7e
6mXWXCjk81Sq263O6mn22SROlLupA8RPVyp/Ag0d8i3GFSVs08Oo0u5hg6xJz9Og
xoEzNOIAA2DUOPXpzed52F6d/Qra2dwPe8FTdiQ2RAJx8R7o7pwBX80Z1X97sPQo
serObndvRBJ5aCDHJdbpaoVL5d83E73DaZlPk5VVOnXsEPRjf+dpYgEV+PRX9/Ps
+7e+kDQ/sJ/Cg2dUGuKzMZN4Q44+ZgQ4LApuWvQtKZpPmNdsSXZfp+9YWCzZPcpd
jXgUycd44FQIsDrqFXu9Jt1NUGCT0hokQ4FXLZXw/kTZfFsHD8WzJcRNEal47CLk
/A83B+RE+7KGfKYEXYRwgE08KGu4BlfyYjysrcnRlbtbk4MTQ5h5vw8dMm6ppZMj
4mH+S3rKBrS7tvqJka0tCazJfOl8rUPMNUGiwzzt6RL1sOIFVFu41UH12QgUGVJy
jmkLS/XDYEUOKINw/S7nyk/XswwA1OwRlZ/x+vgjaCzkmnZwLTjOxtmPFArKFwbC
w4CBfu+ltKD6Wq8x6ZQN2+WD6RTEBk7KW4rEBsu1/3Ho4VQqxjz60lvmdHFaSsiG
yZZMMhN+56MqV8WW2WXWdxezcINNSSNQ0n7LEZ8/kzCc/kfbaKJKvdcr//2w+qcy
Zjp2MmwwsPdksFTYDpsgA404l/Qy7xbf/8CIN1h8V8NPLdbS2/TFeMR7zvLhhchn
0sYhD1ZU51eZhUpUmwnqCjE2aNeLk2LIudNNHRJlYgas1Tds+BubJyO2dMdPnz6f
XbthJJwXxKI09kgKfqaE5qmcoVL/mpuA5XG4EKzqjiaQ/XJysiNuB3TaGT9gHmxC
zUGdDN4IQ4cLKFR6PVjRWUs5jJfQFHPin2Wpz3jOGhKzq/JvXwBRXV9jBPfxdlid
Pal+9HbK4+LTbkaXY9YtxVH7eDZDpS1Rjllr+1gZK5ZOcsbxaxlCk/XhPrEYWw1p
6YgJNfA+B7vEbK4yi+4aak/nl9LQZD8AEPGT3EUGDC1GD4m41I4eUm2IGxp6ye6+
4tyPEODuWdKftUsZNALf/UfUD/qN/KA14OGnwETKeQ5ieCxOgkldrXFOfo0K9Nfi
ax1iMTRaQ3MAMNhgnZwfjhe9vrqKFCyZoUH8ScEGMmoCB04jHlhcWk9KshRbD5QZ
vtmN1QxsXSsoMwZGVpZ+2xPRuRM1ec2k6+AXvaTdIV3u6EPFJo0SYmk9FPqhAbdv
d08DLE6KEhwgljeTjvHvdk9FNAM+I31VdgfCIhXrIyf5CMl0vOwc0nas/CFyOpkm
7Z/ZPgDkPywgDuj9iZDiIDzFTlvZlt+d8eYuDeQn0NqHo+gylfX9PHe7XRJBjE24
Pjr9OMkVVDYy7ReL+5P+v4W5CcTuIXETo/zlSdKbSIInbcKYRTiGmGdQe3IywqN1
alAd1u2Vc/Ls25eKEk9JRBhfbozAhjzvwVZ1yft4AnZMZgWxCKeh54JI8nRMR5Zv
sffHubC3RQ6TV9YeODilQtWPIHOGT4BRV9Ya2pGJ3dqPCnjRrlaDbmSjgOQReBgl
HsmG4vV9GlEEz74Ra/mX33+y09dZGMMGc2qtdjAL13UxgjuHwAL5eQN4KmwQQS56
pmdI1DY0mLwPECeaASNUj/Q1jYOomq76jBw1KUeBfn6MSM+aTOeK9vSaCBOrrlH8
4Je8fD3dZPmL3BoziRHDSVeYRDWw0pUK+w6S97vyppS1LBu30mz305o1Is5ZnKk8
7y6aKCMfnBdM8jSLJowVzBY0QoQ2hyjyAPPNMzY0H7pFT4oPsCgHlUICzKvsmX+A
ghBZ2iO67lezDczI5kE7D7Z+Ake/F2V/hw9x40Hf2FQGo3KtfwdCWUGQhRNAHXFi
pfBDeSDnrKtMNSOu3GGl+9s7E7s1LFvIiCeMDK18lR5cF13AoV8nh8GHBTnZ87YP
KA3g++6Jtk/ESXPj1U4NmJnOMJCts+u5IIsNy6x6RpSuyR50k8lQKNnsbjeFABnP
YJC3z7GwQZ1utlDuhJ4ZghY81g78/ihJlpJGZBElWd2u96kjgMfv0pap9z8o/yi8
x6yBtSvM/zwMZVRJIwtkL7bb+YAgLbC0vznpykn5afwCHFyeRbAa2gRCOAVGVD1i
TagsdNiiC7+pa6O5vyB9uQeXn6QNMpn417mq/yIOgFK+/llOUmnZYZl2Vz6L5sW3
fdJNv4upS3pW5cLXKYOdv9Z59T4E+fJCYzsDihThzgAJzuY8rs8/zdBPdax8P1hm
qy+ccu9rKdFG5vPfM8I76lMHNeNvUbp+EX3oU5Wt4AoSmkCq1+gbiXsZ5EmtfOY1
weceiHLfoTImMuUwLGXgF8rYG1X5iNqniFR9kAKDPLy2OgtqO/g6L3mZnBoe1u08
KrazjY5agYfNq2O1Wk5m/GyhixXZg0OYmCETz98dFyNiwNCd0vRE/ZpGmQLdym1D
niLJakH00x/8EHuilBTaZtuLMrHlg0IIfu+X7E0+0aEQY+os1p3VAjcK/O29suBV
8Ary0ioA5oqjcdFLgZMS3rpDKZeig78yB8zAL0/lGfGZ0YuMYesR54AoRU73X1Sy
SkqSIddV1uTo87JfRf0GvbDdqdtXS96XDVyRlb0NN1ddeRRk2oYfstfECtepfAOj
K680fF6D20CVbEhsIT0l99ptQ0zEY1tEPt8A+gr4sZjPsMnzGb7OK/JJtg29AlJi
yYv7EU7sbJvM2WKVWdvOFalazzyWh8c+T6q4kk0u3aQGHjZh4j15WekPwRSv8xbI
cPL2UYxoe63bCSkX3F/ImLySFa6J3+TN6B8/CH2x8rdrp2v3CGlddlg0toeYekLL
n2loC8SGcgPhNWZkwCi/m1S1R+lIvlQKJQflfwPmOuxuHkVP9pykcblvAUZwofEg
7A1kJtXdXb8GqCPrZBetjVKS2yJNTndbXkLqMnEHh4jaTLGI9bZBcx3Nn5E8B7eV
cxeOF43UPfrwedcceL/MOdNA2JVzVY/FChZR3ccUeS2fyW9eijV90yAqc7ownC0Z
+E2xdeknvNcDzEL/T7PrTDHyyYJynayR/lRIiwrcC+zmGagJlpvoM2hYoZDKi2LV
GvRKbqmCtcclcDa5PqdJ/B9JsKrdqWdIEdMkzhIvFU9ase8dc2aMazttwIPzSMlS
lhqQp1EtZf4joYYIdHoSn7YjD6LlqQEj9dCc8TKxdRh1OwdrhOvQtfpLF4/bLYDZ
AJehN0NPaq/QpyzOLdayuKz2gyvwa2esECJkJkDeuXDvfNUj5vOERBjSdiufWqNI
tlW7aaWxw/tC23NJVvwYix1e7LoQqs/gZ6SxD3MFLjgiyhpu2XfU0BD/D2pwIUo0
f5TGEqN5jzZP2lBgo/lVUY+d1yhd8T7hz3xi6oxoh9a6yknIqu1gG0wH0gOckrlp
5gN1XfNcqW7FejWf7sbAHCsQmbx8MlmRNm3q24mjsOa+4r4ghJ7MWmPpNBb3/aJE
o3iW5MkWango6FFU8l8oD4HAbkGCJI1Vb4A5ONbZvhC2RZVEcPJMoqo2DozS4Y00
jMxQMjoqlPNBNmDaxTbDZPPsyV01Qpvehv8C+eWdbi/9P01D6YV+dIRUlOuZEvul
ez5Dj40iqLJJfgeFFjQhywZpd1JjHZSWATl3SX63evhJ7i3gQNn6A1bfd6P7y97o
0MvFen9Uxh7gkkG432tP+kJqCAtEG38czWj4wjiJwR6upP102ycCnfQCWCl4ujl8
9QeEXOB1okV6AKLh2Ty0vCUWmLlxZdrqCdHQLGQB+eodcih6VJmWq/QKnz+6K/cc
u9pqIkgtAvjeViTS+p9K8KCLChY6YPwO9LtQgIR1JJqO9dgWJv+zdMp823J1ak7z
Zdav4MbNIVPUV/ch+wX7wG7G1WdUexFjMcRsaj6GcwAmXwOIDPEwG0UVC+Nk6mGv
QluhfbjpgX74c2QOitFVl2bE+Z2noPwkX0XboAQV8cOdQko5ZkpDIY5mx81yh+l3
/nRS4F4tdQRLdg6nKwGWPEptbWsY8fsuggWYlvV9RTHI/S1Aj4Y/sZYsVH5+UtSr
8DS5d7XdYAiwa18MC0ZixEl77LyDXdK4sZ2j0EvjJO3ntL6czzmHmidyYA3sCv5C
l1pdTPwtQDA5xu1D6P9ogZVWjrgmo2sIsBMwzkp2QFQ6QkKISf18s1hqKtZIVIr/
SDTj2WV28WGuXjWmPTgHoIPkde3EaVBeuYVaWtKzNQX1jGqw/O1IsFGEKinA+SLn
9uPpA/YAzULfjglK/5CsLWij/VWuLgO8WxMTxmQXWcBXFrLmNpNvtq7WLY9JtlRD
Nn/+ZeotZET5JQ33fsOlv2MGQm1qxo7Z5gkdDVqOByufe/RDWJmuyn9VDG2uSc5x
pR++NQF1Vjt0j/fq60Uq410Is4p7AwO9buDT1/vzihvQKXObXsUMBck278zhlHlP
mQ+NgMYcQjXr4VnzXN8EGCVtRhIYpa+V5CcBqWqx/9Jx5hZNVf2EFKuaXGnGTpEs
femDhiSi1IF3Oks6ZrlnqPgoBDU5SbxM73pD7umEcwSW4sKWF/sFCzLJG+SngwwP
kke82O7pE9G8360vWT5fmCzZY/EyP/tgUZ5ITLkhcPgn6FS5sRRSZ83z+lApgoqF
zXGfQD2Zp53FW2DrWDvwURvV9NL6B7qRgrAnwKYMBne5R4zUb6zrxSMlsAwPfVY0
Ndcq2Ao9W5bVYyoDwBDTRwqF1M/HRcQz8b9yIdzv+WGrdgmZGgWePQYKtY4Jkwtt
xmrHr2h7di/579iVqdcZ5GYkSwdTLfyZd5uz5XB6sholHm6G0rijFg+clk6PAJWS
ZXObqT8r6JM3h/lQbQEUDJLiI0IYe9NU0yNjeYbRV5scWSAG2afKCNujZ+vpkcMh
26//grm+FxKPppy8/CUryCEm+0HpbRxdCfmUFU/L8bRpHvsAZN+6EmHRlZv4yfm0
O/L3NVV8FhB6bSukg9H9vDoOdmBXEiBDc24Ujf3prct6itPhYp+JNga3iuCDNHI4
mqSXczGL/UGyRdHVFUMvuoDCCcEKYcLm8COfIFT7u4Fligd/52/RiEPmeVZle5QZ
jpzup4942rz+7OwkNe2bgdR3/AxEitNrA593JLDhkyUEqNn+XCk+yruUky1AUxMp
716jUR3d73Xc1I6a7aYjjBPmqrtEdpQAcDS/LUalLdgId5CQEIoYDufvnx+I9GA5
465CYCYEPTY0Uqm0UKeoqzBffQvVgX/712ZhswuJg1cuyPNYnmT4Pdagw3ryoJaN
mGKfumk0dxexgEzlN0zC6sVdgeeOMWTYt26gP3JYfvJ9143PZlouSD3wVbD/BpAw
eul1lo4AoZ45HlVC8HDfoexj93K7ANJ0LnYeuMsoyhP8Wv7m/zGLol1NBgjBDzzg
MAHlYz6DOa1BWvvWtOucuqt0hh5bvaeyxyR2dFSzlNaZRDvU6ZmQYSy2xVhya+Mw
cDumziwA1qQ2OClB/KkiDh85eUkeJvfDJ6brikzGXEyN87vSIspKyxk+IIlaedvp
Yd+z7jhOeIZphFMtDfFeJG5kYQKDV3Hd2MqFwQ6XXTprofwjIBosPQj+jFxu4T/Q
/XbMKnBpROS0epjENL4rcB2Lv7otjSoIfp6m/qCuoNsQNzLQIMnf0oYU77Tja8TA
nMNzokX4itIoNu9u2CO0kwUtiK6BQtuezCBGsQSsoYS0bgeNawDNuvTeTyxk4VGw
saERIybQDDYsjMnXnAUIxOxz3nUrnozBtgp6ZH0hlYmDWy9SUjQfpMoRseKzwxzC
Jcu1HRp0qePAZ89OnXd7MGzZnsJOkz36r5pTQ5hH6HnJRUBXIxe4JYK4NTMTBVzS
W0q4ldzW+jEVlcAZbaygsqvjxtlEoqLi4yXt861ZXs9ADUoTeVWjH4IsH9Vudtn9
doM2AdxVb+D9tT7O/F1SBri156X9ZejpIy47I+QUWqHtXGAqsgeAe/HRHstx1h4y
BlyJEAmm56tV+XBo5xZKBS0karvaKQ9F923nWgeZPLeU6nrlSAnBhPVqzcKI66+Y
CSsw2xIUNRDAQ6D2gPK2qjObn56RWZGsbc4XhjNF65mu1ZmSSgTXcSTdoUKAz6Uf
BFotaDYfk1bZGpp8LgNToIBK8n+Zywl6aj/DhhttYewecu87ewNPiZkHhh/kYzMq
jL7X+cJ9FOz8QBp52av36lMzjLzj4vRyi3VuWjNkciGglMaGTlqRsUhA5W9wC9zC
f4ljFIJlTpsLRzhomP94PnSGU5j0yG1USbYsWmONrD1FwrQX7X/i/VnwXDmVX+Xp
yDCLHTmePjfRzBSBeYmF5rxCueAbvp14k7qK3Xz8MiC+kvgwQ/FlLTQ7MQBn/PNw
8i8ZVx7GqZBBNklgBUlZRQKzjqSHtq2QTS4EVnVdErUqhTY5qFmRc1NC7PxRe2UU
kHUOohQZDFpAtw+1VJxbk3wGzFKUMBbGeNksatFYt5uyk6QMyeKsGLiqVottRQbN
WSl+mJ7TdEKVlQ2+9Pay1bPMGq+Ykq9JkLuIsFqRUSAoBQMgz79ALOWykT3Mlqhh
X+TgUkfNPNedyYImR7onbyoz/yzLBOWfi5+OTQGosx7JFbgeOv08lBQVlmUsfqNZ
IjaSZNor3hKLqGldP4QHeDU2hAHSwYIvx4E+ajoAIOeypesH3G/BOFLSKVAbbqZ7
n2eXVGrHWdEFKjmIBaD4s74OKaX2m6G8Vhz+cFsCPgTtFt81MRo9fgH5SndX2lHK
DGQzopTnTnC6r32tT0WLa6gqwBVnDnpwldZC3lV+eiFqwRXA9Rl70pMDYzmhw3fD
/IjrU6a9Ir4tJ/W7R+Mor9OmNBRXrR7Y6UD4QvWYeoE+TTgdLmIRmrjVP1mpprrR
hffjAe8pTLNG36kHPvvs914VmaVyYiYs3RF1rDm3s4WLRTSDnxH98rWZizdD2suK
OpzVaMCHBlFY74WIYSyrnSCcOMB6L04GiPkC3Rlv4926kzHtcUGlGgG65EpGvzp5
Xcy8YmjxZ04AGu+FS8YHy6vKEF1HAiiD3M3IQ6VPQwllU5uTv/w+hNO4YYgqMvva
1L074D6M+aEW+k9I2suXXa89KLCwbudbhIbwBRlwIYic5UeTI45FAM7Nnk8gymiQ
sEJ40Ydp1zF4S0zCwwmct7z+XSjjqFd3AdAUtXmPuUU/MypFMuuktXwc9MKrllz2
97WNfkQCWS+gKPz17mdPlNol4tM7kUUabxdDCrqMOi5lJ6NtjYa9Gmsn7BqC5Bws
bF1n5Vkx2pdawfn2mV5SNSv8UaX4ziWl5MRUmQk78l/BtJSS4M3ieTgRVUP+68lJ
Ih/f3ocEIXwkM3oLwIVglSNzYEzGND78yk4oICdLeVcHbO/2bBJqV4DyW3hU0sCj
hLfHH/cZFtJ4KlbjuVQklEp/hfdme9TsIEftqaP9kBGCAg8H+Szsk/WZ52P+2BcZ
58F/h4cbu+QayftdTY0tOMjQQL6l+XLrvASs9MCuQaIJwfIi8wcJ9aLzIxnFVm2i
o1UT+0FA9sc5lQ/CM3WdbS/9GgZ6EO6DepS/tdM1wNMPV71yiMGOkalJZao+C1x5
5FBBaBhBv5D+OHjjPYkVMje/8HuY35axRv+EKe4ruNSXD3wncpQYUmK6YYzxdkh4
lfk8q1FO3U4IzhbU/SqkfeNlqPhEx9031bksLGWOoHofjkew6nPb4G+VRClUnNNG
xLpQpQgqFQEDhZlNxt5ZZ2Ber/ToMc6L1zWOewp/q8aiFZmcSKo/w3JWCNF3fnWb
jXrDhaUODD8ShmJu6PFV3Gco0SxWYpGBkcfYWQSyXbBunkKVMudps2RlqUfPxGFX
lEVsPLGapmRx1hUKQRHLT15GblSuDbCHrVHWcQa6a9B8odrDNsgELqbs9OVRcwVI
raGCWVXXXCYE2Eu+DGZ1oILYZPcFlEouvMr8/uJiHQ5mx1kKuaF4gKKGXVFHELrg
Ho1UuFp4SSDuBemn1VtBtmszeFHhlMDD1WwM+0pl0U78oeyK9GyLNZxz0M08RDDI
SbpN9jeGq/HtUJ78gU3Qu9zQ8GODK1XJtnV/H3KEaRiLYFYQM3TSg+Ggq2GfZaso
MWs2KQZHGQ7HvX5oKKVu49CsqSlMH8I7vA36/YNyC6fXfkFF3IK3WPvYSJgvOVS8
YlbNJujdKY3TK5vR0Kvz0tu3EitxM85oB971VP/faDRghlwpdj0I7QAj+w5fXI+5
t+kspAuKLfIdeV5jwV96b/RndZebHGMo+hU5hGOD7J8oXhotnk8RgaYvQM4gnUSA
Mt4xE9Kr4Axj0lH8ldCt9gqqX7298Cg+0VCaNZac3DKxCiwxjuuEUZV0KRyboR0u
geJbbpT9k1I7gEdDbwDUPIOJLCrIQ411ZlqwD7tzCFyudvtwA4PqxOEz6KrCaR1x
+1L1IoAnFOAPpdUj8sruPC/zxpCrAFRdMlRxIYPIKc28/1KaKAmeSuSx9YLaEqeN
Mam1DjQYyFQOp225Xhus27VWqMDGeiAzkzbPdY2YT0vICVjNigv4fOOhJebjYQl5
JGMTqHxDgWZgj5DREgZUQWPCAPbswNms+dFHkRlXySxQ0M9WnCGq7989okqvlcII
g+XvONU0fjkSw3fn/IUY3uM1tlhQmgD9NNl8ZiwSbJk0lRxdHBYNWhfjl+mxypUa
Cb4O+ukUoYTv3qFpC734NzHvFIjDda+j1WHxpjrAEITvbviaXbk27v31fkuJ31ku
aGpqSZdfmmvYsKs4q6Ly5LWQvaRwDkDNdO6W1O0TNj73CAlfI3W71wExKFtGmNtM
MTfJABPmQ4WM1yNxs7B5QSFzKPUylk6kB8fATXDxpuv/WqVNE/TN5L/08SswljxG
VaS5aQylgNM3KNFeWiE3I1CIyOjEK3m0EItx2X6jkY3So5dnWdZbcHHY+5BgF5u+
qtSFc3WGNLEdXlk+0IACy+JIWDzoXaGF6wLYVedG7Esau0Yc2evMvqd3Qr8JOs5C
zAqpZJGjNI6gc2IENn4kn2fcw77GGH6sg9UmC9w5aXUx+bjbfsxW/m5qOYANX/L4
T1rWrTuesRKUmkHRZSUbYLKyZse7LW8L1S2UftksjtV84L3DzVxwTnqrzGxtj1wE
9VpuQ0tzfl3iOQ8C1BGGro5N6we+zrBRvV4GexYIf8y7l4olpLLJF2UB70IJR8DB
efKXQB+AFJzthynCHObbT69GunOB/RyFhJrHvQYPrbCd5CVN6lqdS48rsWLl+lQj
An8JMMwh0SronaJPPVAQGJtY4MRtYmcM6A27cuhPySYWWK4ewWtV4lX2enmfZthn
hiDxksT5hZZhg1+zeWuiRgjXrVIE5kuS3EBMTujOY0noFnlPYviP7RnKfrYfmIDP
qCV8sHxpJLSnFpli4dQfHGvz34bbZNAty5Q/o4OUaxIbcYkbm8hT7oGvar5YRhMR
Fc1kKl5Zgoh8fbwTpTXG9tTMndgIOHXBts/cfJTNqiJ+GadfnmmPiexz9q93gmsG
ja7eB8hKrUVIPNkhfkZIuDtER1V6aBWqa+pPB6A7nxkIuK2NP7dsdUkOnM7jqQKM
ZYgSI4Rd459JSWSdQXLMkt2Gu5ar+ZcqK4E6SKCLJXMlpvRnWSOB9MAZa5HfFezb
su3gpI4tmDUfl1jyz5N77YTFk8DFV98FW9fmfhrxTTPpJvFXzvvz0xj18iLXhyvD
uMegq0oleS5pLDX/2F/I/OqBuDqED7cAwv2ezdHwr9P+9qqHOMgEua5YT2bPD5pc
LaPatnQX1z0cNAGR/gHD9kSPfkaqacgrbZM31MrmJ3m0tu41iA2FR74AAqei/cud
4PmQO74EOKnReZ0HI0oDTq+as94C3yaS3Ks+MjiEcGDqD7h2BFFxhbTb0HOaJaWt
HTWqT4nIedLKaQZ0P28qWjllb2XYUuL9SFkOzWQhIhdx9ynitLUBaq3AIX1lUGaj
vaVFfpVHf9ahl2ZV5UuIFh09pGMU+yGDau1j6GDy5MJzU76MNDk5rq9zLB2Cro/P
KQQTXC7jusJG5afjoe9WH4QD6wAyDuOrujz+RJ/YupJn6vqP+ETz9UCJGaMeQHIm
WMIoLTCd7gtpTn9rKyOWa8tkctfo5IJ9GOa8b2Pw2RQ2BDSx60liHmJjZuRkO7ie
oqgY5+895Lo4iHGrw/mhlgnEshgOYAOV4kxWkCKI7K6jB8lzDr1NYBnoB1L9wR+y
+8QfHal9qEp1ClWhYI2sKOH57vBcIbwf/+npn612kQ4ZiCJRcDREUcM+JINVkiq2
m4OPuxqE1idEWzBiUm140cLWeXGY7n84d6vcvEfYGCRTfYYVUkA3r3S109hC3uie
xO1is4OeAws8CF9sSTNnUMQ+f3dEzbubrHyWAd2bz9VcQkACOlt9nY731G1HANtl
mYluSExqUWRZ8Jnaq9Jko/dCYi5OrRC9FbU3yWwl9u8Rcdzb7ZYlxmUI2g0MDOc0
dWOclSJKRAlKHqzIujvdIUmbQSPYbu+ancM79TycKAmg9Y9e304FjkGRzYqR7ffX
lkMWq3j8eU4mqRARMwiu4bQ/nuEROQ2BDyOtDK4LPQreX+tJb4QFEqa080yI5ouv
d3bHrb2XRn/5XbT++KeR1/t8xl/6j8/jZxnpvoqetfReIkOXpSZYoJMxuVTd4f0q
tNSMRybTqWbS3jwx3AYgUunwa7wTCTiTojMQ7kXt4Vz7R5BrXLP0tuFgfFTskDwQ
JQKIqakolGo7CfahAafiBlvztwizPcFKHiHBIpYrutLcUj5WOMWMdVLMx7z5a2+V
TmusrsjF86vRLrbXE1Knc9vFjPJvlT9c1ShV9vhaN9yxmIyKtlr6iMFPqfGkHD5+
OHumLAywxs6shqAE92Yex77o7cUa6HrWSpGPJrBZ0+31bJVQLLpeOFtrZYloYQSC
oo/G0gIesSbHwWb9bKfLfYH7evZWvKt+LOINr3Z48EQDoHovBJmxqO8XZTTRSg8z
aRuWH11/+yAtuYdv1MWwy5PsLZ773giO5ukqMiFStIfDVcFe+BC30HjcD3w+rPRN
k7uDa05G7NVOjy07gRBYKZvqAwctiM6SP6XqcK03rH6/Rte0hm6QyQosxFy1/3GA
VlH6kiYF4j4O/MOYdJrWkQ6B30ObuX6dvvuw4bRO/OIdOfSTE2yJN7CSa1c/8Du8
3gXFE/ntE8975ZsR1olf+1BRbvdQqIEoQZA6td2XtZqpnH4yvtaLWbXTyhtZzy5n
Aj7siKlXC3daMA4iuuOYKo0I3CCRTizjnXS3Gj2rUO68WSv9y1g2m7SknKp1BZuj
iX2CkKBJOp25tqGEMLdja4qSIHhZO8VceDEOcqoaYkMlOxDaTuC1e/3WQCZGtADy
BlhGaCfZMQTtFMRRxbjk10OCN919tZQ+0KrODnEFTEIeWwdRUlIrsz52cOEbHhpD
sSVoUHb7MOf9BJ0qeazrzvqfxv4EvN+r71N5j34L3GoplODjnLTAMCF43P1wauWW
+ljDnkNgIeT7DndwQ8oemk4rAOXXwgng23QKMtSAU70+0T6ngY98DIenvY73Nkg8
x48x1k1Hxs0+gU+6gaP/n2fTCpBohZrlUC8WI67UQihbp7nIm27XZezhqOs5XCRm
Bienc1hhFxYyZwOCJXpsD846ZaKr+vHCDSIWVuL3XmBGo99OK0sFBJ/K7VgKHfx6
Ar1FN889ABPRVmvRo8/xgEWgM6I/qZ61KRnrZeLHvFrJ0mM7CBCCU1Z9in1oD1IR
NTXFcvo/kyY65RnyE1RFisqzK8orr1ERcp3uW61EO9FBxoyA4i3Iu2xhzo3c9jBu
IWQHOHKgmh0Dzp2hhIZJBLF+L4oFOp3W4HQmlnvGo+NsxPhjsz+H22Bme1JgPmdt
xF8WewM2pa9R/0Me1yzkWRA6JCIOWQbwmXowYO6hGqXWafANAUvsm2+yoLFdpVrs
iioxnriD/VggiAG10ESQtpMeyuTniUxPDRY5SWu1TBHFELheW6gHe4UnjPVhuLZz
zn0Kca0LWxD1RpGS+1GUAoXFqOdBkViHb1yv5GsXfombkfRbjNBvCMMIRQZaDmgL
9iVZfP5pS4+q/iqomEnpFRjphX0Ks0nKEnJZ6yFPEKfhXWsqXP1ZuN6iLGpHbMkx
xUOHb77gJyfxEyAdTFMIG0Km5UG3d4E0w6To+rkjA4MGYN77sh1cE601M6c5wkJO
fb2JKMsGMOSIg9Tv/br10W5tQbDThVcuakX+UbbzvOBWb6ZCXsyV+78cYVr2M2LJ
6CAcUZ7a5osKrMRvZW2Ot6lb30dyEYJBqrzgoWRhQErSBEeZZq03XusIggOadTyR
3+/v29VNP1ZD2YiLMkX5AounkulvIM/Cv0gTxVMm9BgBT8+OWluCeecagp++UMrQ
th8YJxNLzLByrlILhI4dwjyQw2mh8S1uozSaLRE+figShFo9Id+Fvyf/IjYN0x2L
D1gxqMU16DVXApYQTkhuC2znAo5BoW3c+9cP7Rt9jaJ25N76TMSM+Ma1dSzkmcgB
XwFW9aCB5Fi1hJ9bgGmbIAmUQizKaj79c5wucWgjWHD7OMvhh+bfKPAgGgMn7Pzt
Ev9kOEgpA0oDWgn9FyJseoij43yUWkW68znE7kXNGpD4tHnEH7ZrD8DuPtgXIA+B
jcksyF5fF5UXylnTc4LhFmn9JXqNSFo88692kzb8//K8qqw1is75bW3kiRleA9/z
lsysEIkXWMOjNx+8Ztp8P5npks2TU9gBgbbag1MhIXTFrtkVPVVUGvdeKe06q70a
I0bTmrDs6VbMn+K2vjV8tyFwUy29j+tdQ0qsv30o7tiEZ0SN7o7RpMVimutWrNiW
dTEeNajY2jWLFHZf+0wHFOPBALgLBhtHY+ypXkWAhsAB5jUZnIQyw35uwK0oaU3x
POH/upgVnPDY59mbQdfhYOFNDAT0a5K7Imv0Y0aou8Jr4oV0L8j/Ry522Yw/OTN2
/5u+LCy5HO/KZT4NBaFH57z0QOb9BbsuxaWvvXGbnOBVryFvjq88s1eqMj5tfu60
gtF+B8wtPUUgcWSMAwUS18S5K0KPb3oOMQBgU7/7c0VOXfBdxjuZ79clGUSnLJBq
3aoTxpVXrWXrhl6+mPUTT2rXJmT9Fm6Mp+SusvGrk4sGxL//uHtRiAbrr3YTMbql
KfUgTW34Nr15em/hKHNYkdbHHZ32VBF5pk2NREy0JMWeYpNx6ocQuM0mLDqB8JGg
L1Fb0yTbLbjj6ohZy6fVwfZ4pcnyWPuj7MvaaQ6KKLeuamJj5ylZEGaJOUJY2jgw
pj7kkAWWeiKaqsIkEJ8dieAza1qKRv5B0O6J7LvxKTDOu2g//kMrFV+Dww6YHBgU
MQ6XE5rNtCgkx/uA/ZKO6EE5cQ79W3iUR2xJd4HmGCvGRDlLGQNtvtRZZCf6imkh
J47YrdJxGO5Xr5M+Y2sebmaGFs44FpD5Tfkp65fahc3lv3o0d27Z5SGhUsnY5dTi
IO/TNFF5rPH7nYByXs996VEp1+lLZYGojwX/IVGHuKFMIxvN6dQnAeVPajZvuTIS
2DGp+wWMOOcLZjsWX9eFYdDWW+eQjcCD0fAwJcAoC7Yrs8wwo9Z0Rm1VeH0kw6Di
4wYhlK8av3Z3+t1pKI7AXlnWZ5gRADMa8F7M3MfRe1XQ8s2E9OfnJ0Vf6TNtw4gZ
aerWwH2/VnecgTJO+tUrCRK41J3jcyhZgVEYuIeSxenhLpqvYObf+gjjd65oJaqF
s0QRd5BI3jd7t55s/VLcji64pyuEVx5hh82GAhoOpX3ddRZg+wDWFDj0i8py4JMl
oB96Aax7q9Q9FVK703zOYadf1yDmgu1lG6J/mr1zCJ/Qsgeqwj35U25oTO7kiD80
9fgLW+zhNVmigQVdmeOkdw0zbIJfimfEGSLvBl5TZ8lhIyqgj4hWjo05ytqsPp9x
v05XSjmdZwFrr2nhuWXMdShqOGeAIgjOH+llFhaA3BxvPSIvDBYGjVTgECgz47RE
oiL1IhfPfVyhVfjuiafQLu4XxzwJ2Y+7s6YW31dokXlXzWW0qT0k8J5wBDqZkiBj
pe/zNIjX4abvzEJAtz0sha8YIKUhEEjpszp2J5kEW4MfzBo+aaw47Cnm0ySoiyRB
TrmPz9DVjapb3tUy77zCGQS0eeBC3ziQAtEoO6Lg4kiESxnQkRkLzbQ3kUyCDtxt
i3f5LDF2zdL7xliUH+UoBO9psQqEqxjw1vRXsS52pyVcdaQkVObuTvvXIy697GAx
99keeeD1bsJCr8HDuC5uy76pMe4me3w98qqRsJaCahJ2Hep0ppO8P339bLUCLZbv
3W9Kfj0sgdfcwrcq2Lhh9w0168pGjC+AV057txhqBL7ImxAYXqL6L0ft7m7hfQVu
mC70HBHH4Y1XOb6TQDeSW3uaAFJHGBuOBJzgSK1qFhC/ajt3U8ZFVWjiPNsl5+2c
0dC2+nFOlMFDRQYW5IPOQ2lXvIATmZi40thHYItM8gc86rqla9NTToY4mFhHY3kF
k5E6rOz2FhBdOnHuURIIubikw0emavH4nUDcDCFve6B6qGZJziPGx1sgEaD69FNM
huxuLyz+pTiNGJSkISEm2xBModrCGGc2ABCzwUhtUAsnL6TmXPxBvpkrqvNdG7of
JXUpV7oYU6/PeEq1A8fKBbuMfiha8NvOHSooJwV6qSlmc2fKj1LyF2tLAnjuFxoC
h3C1g0rmn8ROH4jBm+GhYU9bmty6vPF8ZZPiZroNw6MeFRG0SpathDai32WROozu
m0BGqQyfwGLipte7XtXRlq+0dJhyF7PlN4BwLIJ9PBuIlzca1pf0a7nttYhVxEFo
mSSHt4MTqWR3gHZJOg5w/3qFp8mWBOkx7JwCpPgaC5886yQj7J6RqpPz+XdH+J6y
tgagFoJNpY3AE6oBoUKpMehuxuAPgs7KugbHpd5Zv622Wh2a1uWdHtsLh2PnmSDG
MpmXPt0UliUZ9xkMgFJGApLyrtR0ZhRNYwrkA2Rgh3lKNxBfOk/aBhUnlbz/o26y
15JRjPFXS7PajY/ygjSRWDB+3/Mpdr3AuQFOarbIGz3kb9xoUDGK1z3cI4sEH358
jBicHzw6YlcruArhmAeW1NoST4CH8cPsZ6fZYY3JWUWyWGYA9oT0jSDUvfdHP0Wm
UKRCIRySX1SKy8joWUjcTbDAFgnxHfhnCkUT46FMLVvGyGVjzbdbvueWI6DYkXSj
Nsm7uBz2tEk9ZytIFL+2hWxbC4bNiHzLNIPv1BSor2FzOYbDg7jTgRXlYPbrtw1H
/WPzmXCzvMepMMoulSCZPVv79f8FidP4FAa47lJXS8mJSM+MMXdwD28tcdcYIeKf
t3tXHCexEvryHqtXcmgnA71/EiKLku0WsBlO/k8q14Txhe18FqRAxp0YpCq8NLII
X9gMDdnD2QxKeCFniVMtUkpU4KvTxDymGjsDG0Fe6LRM7EA1Jg2z72iFF6KYjE5y
W5An8/6RyFFpKbqIfxPY418wJrrL9Dlvz+7MujPJAn4YNh2Du69vMXx4tlYRLL+C
OSZ40xzZvBwjmRnuboaWYb0pAS/j47tXQzYDn86I0GdePwP3X0riJiV5DZWtzDWR
ohjAEOQ0pS/eD63dOwaC76KaqL3/dN4BCwD6UVZCjFYNGxqMbor7dZeIOtDkOw3h
CMwYhFJxKqd0ePqLdenioTXxNT3f9LTAL1qEQStPJ1P+6nROeHErpDuVhrAuC9ae
hJkO1t5oBYjzXPAbGZ+d4TIV0N2q9DOcoltS0DWr/13uQsObb422bsUlc/4gASAX
1jEN356K/gHp0eQi9c85FG2BnKgm+aeMOHY3zJdDq9vy07SZiInMNcTY2llAN2iR
8CXDSNZcm62U1O4E/RYitvYFYw1KN7tmfyFUVccNHzRgZhleM3TgzKuf/usjRHnK
oicuFfRrZn9LDLkyyZqF88Jnai71x+1nHpLBwa5LPGDSleXhDXOeK/Nbq7VY/Cy3
mcpxbbpJVx2pv3mgL6tmXKy/UPkw995mUL/5zwgWUbD3nW3iBDyfMpjMiM+s42I1
BGYL+Hc9SUXH9qce7FP1FZ4MBqUuXNG4BI36gM1lj0H8IKqFFl0n9umKCQbUnBib
YuANY+FDA7F4KfR0pWJlwa/+beLqM9/jFCWng4FGUMA1Y9dyLFfAJWmS9fM3w1Dz
zJleByqM3vC06GmZLflemidTANvZhHpg2lzByl0xywkc68LuPy4hmLfAWjhCLvrw
UasiMQ2s3YqOsNIibboJG6pTyXv0IHdQXtBXNm35dV3+DaEAlSm4j01SOY8QbIc+
1CgzhFfKyydQbao8fMpfK9pw94aNQAxpWhMIYrHYUebibJpFVbSPiwMAeBosTQWb
zPuhRJ82RK0lgpBllEu2G92UoQPT24BO3fVnm7J7jtkzLodAlE/V+CgcWJSPUQEP
KxC5Eo6Gheb5JXKCWJjR4BiHSShDyZ4iu368v2EyzWoRIsh9begJdxr91z2DCy7X
BiBIw5A86xbnFQubLiVXy5gWE+OZ5wW1RFii3Typ11l4HwEGe7/WLAerWvzep5CP
91oYxjXffjGtnrX5g2V768WpTDTS683RV6ARoJkN88N68Kry1q7VJp/E3eeTin3r
d/aj70s9j7b3Dj+nxpoK8VaskMP1RaOtB8pm9ImHYa4QVDhYp6apKnvwNvwffX5C
5ezcmFK9wfNiRGb4Sboz2QSmSxuSPf/YWEGNMeHEYU1v6HI7DWC0E3BWj9oBX58/
N0Vqkc9zWgQ5lIfCg0noX+qb49A/7hEmGSP+2Y3AB60+tS7gx0W4YH4Ym6kBMwr8
2zaHeM6bch2cmP2Bu3SmoWR9FjGkUhfrB0dg3/0eRnevkavrFckCXHnsESH3N/N5
B+FOS9LuqSJAcTTPtrm1ARUe6QfNAVghc/7b0ZiFoQzbDROE1u8Jrk1+BEPpAh0u
cmK7uzLOEvqFPFxwDhA6xkWCj4C3Ykm8bUm9HWkEgFS+BQ/eeEm+pVE6FmTUn+Xp
QS1EJEs+ymmVIOiZyDfA4adE9Eaxg3LbMM+8YVyihycpXPhRc0RmPtABHUMtCYCY
zIDuYLqRFXjS4K/y6Dk7uLjH4eZAe4bBUGIu1dmld5toWDxS7z0X+qo8RIcIVfDI
6vdpHU/KUDF7Sm3QYoY3DxY6MWOxEDPEB582inayH7kESeNMWIK03/sG9pYRdCil
fUmoNfoE+W+NxVHbdSvnc23OcLbfU206UYMW7+4U2iCXf40vHTNcy67+yHOCqJm8
z4CYV0wPpzPAEGcfGGCNwaNAZGTYObPU1hM69i3CODWcHN/gmeMD6L7UN3wppDmO
TemLi5k3LQFnjYftlHE7o3qU3mnHMeMprZBRp+uQvuov9FhXEzfk5x1dPrBLeBHh
ZOpIB3ZcPtNZFrzdCNvQ8DUT5GlC1qYuwNQzkAiF1xRJ+zCxtq2jGyJXqKPyaK7N
uAGXU15ynTsLTsApSSqoTEQyqON8f/frdRlLIue3dRN/jBW139eUV36HTmN9BfVN
xK2TvVlxxy9hYAqwwPxKX02Ybjxeo8sLVoGnOuUGsBrERBrOXRVRM6jd3oThHyEQ
S/9F769Us/okq8XlCZcCfI2X5tvNZnlTIxEJVFIq0C5TKrgKGgfO5RkXnamMgHM2
5AOc8djJX4lwXXxHBndz98TtPjhgBLuuZwRsbjYddvBMYKXiIjMpFsYexOUexWoz
EPkmvYJakwELsdiuBQ444JL+PRWDCsoxdnfZfzvv5maiWWW4X8EDBleAZuwbM8ma
5gKBgxgDQDY/5OmdnXYu9RD1p10suWelyLWeNc9BCwCWXKXB1woWmZKQfWtcRj+Z
UmsAroisqUY0mWHha0TFPK16osFW09cD+gE6y9mKMKklHB+Yzf8ukolyTCpU2DCc
RczR69lQ/qMCLfCtSQdUEoKE0XyvQ2rnQGLt5NZKnOGI3R1thyWfJty0Ks/VuKMG
zMdgY8oE9HDgYDmjI1uyADCB2a+zbfOZVlfjVrry3leB3K+zeks5W0BsqS3TRTQN
ejNcVDfEOQ7JnlFDOidBU3jqCdfy4hS5igqX/uE3nBnR8vtr3ao5uUp2OTWCOoDt
P6MgbK9WFFGMq72VdAaO/8acogAX5uCDmo9dDK5bYtb6l28/p+SPS5XZNXqnYtze
JK571FYYL+lyWz1P05zHrdUvFY2bKIKwl7eb6UpXWBqQyJNn8xndBZmTQQvhh7Zi
zwYzHI7VEXIBQb/zmS8FgB6/5/NAovI5IX10PpihqfL9hTWJGcje+OVq8aVyve7d
wgVXLc/VeqdgcHsGfqq/pxUmHPWWghFEcA4vx15Pznvdg1C9hyFGZntRGPp7J0uB
ucYmloCQOZVWbxnMICCBakyRLLhk8ca+y+5afrN1eDYmjOZsHGPwgWUe6JLUaMpS
yjiGF8/HDl77tv9bNCNEWXqDtI2YD8+76PJvj/z1el7nmbEvAgsga6QCb7JaJrCo
y2tC2NC0WCWCwd+QlxiSAsAgf8u8xoLUW/GvMkq3LQmopTMJkIT7ntJ7AWwxrYrQ
WrtiOavp06UJJ7CEud2qgV8mqTno2m2lBi9nxzUIcC8V3IHitA21WNjYJ2co+Iyd
JHwglPo3MoCQyQlaXRMyB9nveAuD5pY0LM1R7hFr6AAPTN5+FXp/yu6Fc1AiegLt
UoCsldy1OfEW6YodY3r1RtJzwtH1zT7Bh8IETqhB+LfP3jmwVCzoq+ZtDZEG26i6
pJvLinjgZ2ZARiXZi+7deL9msuUVALhVKmyyM6kTdSkvQQxugQ/ZKtw7hFYn+Qdr
9DTHaR3EXE2V9aTzYbJsbFH8Btt3m2JcgFfyS7W4H2FqNInIpwaH/VSVRQbTDecs
xiUd2LfNJOAJ2DTzWiGZdmPaJkkp/I8xFKXdPOwbmQduid8muFiGNnGdgTUHUdHr
ZA5Qi+AnkixTRI7hthEqOriSBlvInClAIC/1xX1pxoU2vSDQO+AIbPMxz8yKLi56
5HS3tIdZXIUNXi9G1gxTDZCGJaSp7kjsEdjksrK6VYyfzclnbbHZ46hoIy5B2Jex
7K6/pebbg+GmF5U+yZSQY65UokuSeFXeTiTSPDOaI2eH2UrsOZ3TnvL9szqw9ee9
F/oB3zmi2VxKYX/DdUu6XrPUoN2lSxPdenpAivz/80f7tcqnItt7X1JLoJZqzNT9
M1c0Snsth3eK4CQQr409wKsbMgC7FngVN+Nq97uzQz4SNibOYfT7RwBod56dnHub
enDVkhm8JR03usL1H6yHZnFwdKXBcsFvfhg237+e8UlfHMz0TMMT0DHbRb14YSv0
q7cDf4lWjExq1RCeZStzdU2OLBitn4nimn9O/1BURlB7RHFLFMhUeub5lr4ACFsW
q8O+MhWvD4se781g3UzYhXm4sz+V9LFRTi/TzBP7PaESW1pwLWbTTJgVQjWxpbyF
6hebvSTgXG8N05zEWigaetVi6WhTnfVGRcYI/VuG86yc+GNIiXgUfNXPIOsfQCS2
nc7UTgAz2warjCoae/R8pfFDW+ehD07u8z9vvcCLb08HH8kahVBPLIPot9AXcBG0
SbrjkeROCXI7Lp4NRq/8zEWeJFnN5j0cWPDC7MlVynKZHwCoqk8J6LeHNF+OnWXg
5MpRyUoO4mu8afEJE8KqG+GR9txpc9czSTT2s6hsFUJQOKuUJrDqiHn1a1chvQZv
QLRl0cAamxLXhBeIB1YR0aQmoVI4mriZ0w/UQPb4IkeyyF1BO/hZjPnAh7nBY2os
JSNLvLyVwf+06vp59rd7a0T/hhbbVigBa3rbk5AXXGgOFoSQnTPidJr/1Z+sEYGH
/H4QK1I3GkLgUJ7tcjOLHSfmH5LzRfhefECnbYcbqdzKrsW/5ltIENrnMQ2L4THe
g/U4z/Ije4e2DXyGMFxQRZHI28zQeObMS/FYfmKWbTimfciAF5BBCkSazQObi0tG
g/D3wW4tpuonXvnTCDLihfk42JSaom0JqGn+VO+SZo8=
`pragma protect end_protected

`endif // `ifndef _VF_AXI_FC_SV_


