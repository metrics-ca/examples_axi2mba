//----------------------------------------------------------------------
/**
 * @file vf_pin_mstr.sv
 * @brief Defines VF Pin master class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_PIN_MSTR_SV_
`define _VF_PIN_MSTR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
FZ81mNB8JDx5PpPc+Z3jDOdT8ja8ce26ZT8LU5F1Ss+oiO2RaZ0yZ7fHaEEqeYXH
Zdu3oMUTfoTsP3hLpJSxlzeal7L3LDgYl0riG7Wmug7AffeVqWNmZgdzDGZeeWpS
16qldpQhOmjZwtc+pmyQ94iNs0flGArHpHRfCtwqNpfXqXKw9wMgYLicIABu2RpE
rogO+/qHMwAOR63HefQI3DmpamSNCNgev40nRAzS95H/EWX+cTKk0Vgi08GJKiY6
xJ8x2ZVOGyvrqvQqu9AI956kOBm8orgqv76YcS6l6kToeSz0R7rCe53fh3sJZpsw
Q3olowmZ498emn42ZYfzeg==
`pragma protect data_block
JSCBtBHSYIXBA8DEfKXJj5C9nX22RS3Tg6+QDTOnx7mFIjABtWr0A8UjAviY7uVm
aZgHdAv4mlJXx23mitQIowsbg4bYSxggnnzEp6CMPAatCi9zotUqDn1Fc/9y5foi
Vdcwg+jyO90cqv+Zv3wJuqyYWeqZV3OOzLSsp779Qv+A24mtguiTR2yAwVe2/igW
dm+wz45AVZ+P/b9+0lc4yZ5OCtR1VD38Z7OGo3PdWd5QQ4vvNB0kK3RnDAZoHg5P
f2hiViq4AoBzdqg5q5INpbb+9GKbUA5+XCQ7FUVlWagXJ+NhLOYMhPb8+E4ZJPu9
hIJUYCsyCFSEzQ01D7vF6+NaqQig+oXpRtccLYwaynBN1SsyTYaEaplj4vdt5NPi
5znzTyvIqTpFZWoAY8UGAavppxytn4nqd42nXMhT4wUCGrUHaZgzsybhpyz30H6D
CmJrtR28aNgjk1tSWo65Il85abYiQBWPi6/riiNtbZtqFKbhwFSrXBiCqMOWR15V
iYr7Eu+Y1484GPE2UYIGWfu0tR+QbYq2i/UMPvZcLxAv9GVY6Q+fo02CE2il5F1G
meSxZvUYJNy2VhqnfFCbDIguM0Y5zosc3luAv3iGicEFD18yyD/Cwso7AJf1V0k0
nOM0KiLSoA2BmoMmvTZqKDS1pot6dY5y42QnursGC8ExebtO11rBLbZnOnr9IjTV
CfQl0ZoYAIkJNcU7xhjOjgTRV5jdkreEnSgqm2IOpvXN34uQb1HxbgINbigejVMp
onKTcAaD2wl+dDg9mUiu9xqsG/QXQRmLozzaDz1sD6nHA46TPEiAHpqfPuGSQGby
/6v9nHPLPyhuiS1X89QLDDi/w5hNFp9XInxfom2Iv0QME+WO34a7U6e5ZF2gzQhq
OpA4sW2TxaaOo1gdnAb7sAzX4/jdE2I+RpyIz6PFn3RxjsQxEVyZO6NGpeamcBP9
yyenabwugNXNu4PHfQKPuqQyFyJGeJaS4MCcb5Vpogz5wzDcsteXd0pIIFh86xGG
UbC7qQY43z2Epj+qw9jlCJrSmBVZqFp5EUoFyZ6fLP47IsviN/q9P9G7nuxXvF7R
nTzEVKla1WgBWg2OLvcoxBx4fwxY43PcqD2rWxF2nHyeGhe7KDcTYu1Z/OZS1QHn
Zzuj/49IMXyNltVq4F2adMQmzLBCY2V2GpV/tpw8dpbAJ4yoYJYoq4V/HtXfPmar
nN4OcBfIe7wAVOqIBYo0OejqygJRKyQ6/Dr49c3xyEIsUS2Mb5kfaQw/t5BJaGgZ
i/YiSk7Up9ArSNabomijcdb6ZwOUm0FotbdgNCMr0smd8eBuWWJvKGcHe9DBh6pS
K7Y6QcBXD//4deqw2qghtyGw1XkFp2QVQ52j/Y2fRSHlEquv1Mg58wVC3JGpn2IY
jFcGezH2r749H50jzJjGKnjhLSDn7ue4yCeAJglKHYbd/GDCzYHdV7qH1mBK/lNk
l+qyou50heJ/v7ty+sU0+2AsTvKcfZ52SY41HRx4vMF/ZQ5RX/tLqSckeV/4Ct3H
FKrEeJwyUvPan1ATod7HWvvXO1/TGJ9JjC/udxTM/m1VneAbSqfGrGb/B5WCOrYN
Erq5Da8LlqG1dh/kGe9pQ1ynZn1wylZ/GuRYH/i2w8GEUhdVYgQUjxrv5x5gN1bM
0V9qZzN+pMiOGNeTi52sa6H+HzUHWEFuyLiRuPMYM8DXSpTltWlH4za0BPKvW98s
IiqQ63UwEpIJ7rnErvQMEYIe/ZbBEc2Akqzari3dC8skln3j5prVU7FW2pKYxJO0
vHFlfbkHtPHELnmZ64EgQF9odcRE+NonD5H298or0QOOaet0qXH96PGeNDV73WmE
Jm4XKddKiGjTRN9CG/diNlkeZiKiy34KsRnt34Eq2+jGJUFOmUSoQULxqDMr5NsX
rHXWgaiG+qto9DG9wsChAz00rwgxvHS5rwoH7O5ZAVrNkz6G1Tg2PkMk4dnTnZj3
AvBHLlOYmvmKxO5PqR81e0lJj7wB/QyETZpfT6WWhnCmS6opXzIDzz8f24NF63S3
Hp8L6nz6dtOfmVlD3p8A4nEe7HCxXOw5v78YNyshdzg7du5xDnPpo82SeNhGBSaX
/mcAjVqP0ddhW+1sI/NQuP00mvLQHjtLzdjCLTCHsZthjv1NKyWRMM//IwGd+JwW
oCytesw44haHO5DFlzdofCwJ/GkR211ihIR1MxROq4WgsWQ8J0iCWfQDlEy9uC0r
OmqdPzzTIRv2AmnfIbKsyq7P39nxg2Qh/otr5Z0w7AXau995aaDa6A+lbAhfg5jr
LwjJPkOWsRwc7Cw5Q0cU5937WlhjSXX3qMKeyB/0xrIhLO0Wrv9VDbg2DmWoOnX6
Bb3eFonR2cBkyNqIpHkWq4eALVam5nHEgpHALQzzz4G7RzlqKu9FLuGgAaNfKG5k
NqBc2jBJu9J3irSrktTCV5aS5dvTmheH3Rfpa5D53Y4rTAEcJTsOM+St256GQUtM
VNOikaiZwlE25o0hBPIsfE7mzQJ+S+L6rGy+7m9xuYCoFCxuRyDcKQm6IP8OZBbH
80IsPlkHns5leVPKzg3jVy3NjFnTk4JsWK11te8Om67mLdPHFQcOhrLCEXM4c0sX
lEUmbrUcCpvx6YLxs7YGaIha9cHCxkgQ5gD9tZ4cQOzr0Wno2QCkIs2YhxcTYnlI
veg5U6H2GufOWgGyAWIM5WtIGM+/T2dpvw2ll0QzZ7hWf/UMgtPCJC2ToUnQeZYk
VWAzKKL5xyyqjdrCjvcPTOsbU6+19jORDVV/LRJka7s6/nEZqfHzlCiyro0qHhVj
48j0U/4fFD+FzDVi2fliscBVTq9YXgjsxVzwm2I3HFsQk6OD3F72jvgoZ6jgwvkH
IK+frVyIHBf3m67RrUcJNXFMmxIfZ1H+wb0iIwTv1qbCRgMF9Kd0LeZnEIoVmrCb
Um4MJp4JYk7gC7zCpGz1H2STNk2pgZWEygcG07reX2wRZb9kq3ZufjpGfxbwMWxA
Znf5NUJdep/0bgjfCsD6dKYRAz57ov+zN4AYuHUgbGYWEmz1gP45KfeWYVK8IRLU
i5X7uCpNvtGush+NvOtqy021hXxYw9HcMLnwZ7yal6gUH35LqS2o/jUp7ElJ1Ffb
cwvSD2DWhfjRfJxrhpRffu552+N+lgJbEF5QZYiIpKQ/WfTEIyO5C22TaPJ1wKLg
y90IBjG+j+T1v1rNo+27zp2UgJEPDK2eJQTUAT4jBfSJreoDwIcGgcmxQZtmVKKj
nUgh+VM1gfpddPVyRFd//KEY8Xw6h0uyF3OMVqR+U+yOk9ZNpoDI40nwu6CUlIDf
WmcO9vYaz/eTIcdwlpuluOWu7aWbjXOfN1YdJjqFfY9G4c19SQmEaNA4SipWZLaG
TBj1+n76S7S923hFDGNk6VqMJwTHhDi0U1jxpRsSouferVl9sCCvmiRIIiyJzfkO
Plq2zzboE6gXPKlsneQcDlXl59x3OTtmvmSTyum+ExKKJqm1EUDTNyLi+WDz4TQg
9pfodM39fO8zfmQhZwgd1o2CAJUJBPlyr3iu+mHZtC/poZYP6jVPKwFF2kalSEcR
PPhBvK6FSwNcjfkDqNUSbu13fN+SZVqW2GKcYnK/U9dBl+zmUuX9zJWAoTsRTFoi
0VA0QUHcEsHDyPmQGFO3XW/ghuAATu6KBU+qFxyDoKG75YOUzB6KR/+ccHg2Sp/u
NH7tdkdYsOLvX+efbFuDG9USWXmQT62DqXin8z9yhME8JxgWK7qFvkiGBRriWPM6
qhel/yn6B4MQVf2g3BvAyvdk47y3AYfihESHo4yvfyIT/wHhdZ2Mi/DZIUiK3pfi
rOO5RB9Dhbm1lRjvzCTj0j4ldZ8HF1bjBUYUWf+vWO9yHet8jP3LC7W+IDblLfE+
s2uGnuVCUiqrBXiY4NnsP+8+4kxNjOyM1YpBdkjNVpp81beUUV0D8HRzdGcsNFa6
GAi7gDNEk5u6NiSgX6qAxCa5+LeIVIEXr2ovb2OMtriu6EhS7VLAeuC2X0oEw3ok
aU/NiGx3IUlBsrVSw4+0v2OR68CFt+hRXWp8eRHY2TDMEDjco16bU4aR2PRlFdWj
IQkWa1LCIyVKyDD9fJ+r8MgyPK9QZbBqKvN3C9uUiSPNQzGcvWNZOa7OcxvpSSxt
5EKxJNNNNeW+wDUrG2mwzdZfHHwMWk/6QLmJ+sj80WkiX0jAyMMOCVQrIy8MX2u6
fc7K2w9Cr1IIp5IksjG5INgTeEO3hzXR0dN2eBamaFow+Alf1rmZ/MTlutQs4YmF
NRab85d4H6X5Lo/kOowb9y3o9dZGAMctSXrjQ0ed+7uzmRfCbt7J8EqZnlK4Vy9F
b9HFQ0T6oEDDI3opvs595ql1H9FUns8o5hds+m7D8VzGs6Su+RekshavzScIB/Gk
nMOT2zylMElFClgq/FaI4jBGa6GLYiXJl3HEVmlRHRF8Z/6b5YT6+fQTDmeZywz5
pSmF0htMjzVLk9eodHtHvS3JG5snOiaw2386n9YvPL7udw9CQRXzeH+uXdjPUVFH
5TLUBglIV/j0m/vhDXITuta7rF0D+fn7oVaIW2mhU70PusLBYczJyEd2dng3yKPl
5pCzSzGoahJd3cdoLY1alwoLYRDP0tu0DkPmq5dOlcWH2tnfhuK9nZyJSo7APsqn
CYQ5KVNCGMRDbzUtqZxp/LzDs/BMc8yCgNAHl8VI62icA29+8vZOjbscTj0OuWPC
NJke9VH+lBqnryE5Lb/Vn2hfgmiRQgCVW3RDtxYQHL6yF2VU5HCMT0CWItdNf4Uq
Bbuobw9Z8aq1n3eJE1O5lXj/UiZbMM6TWs5E5/6QCSQ1KdItR3a9eGLyLMAGn+wm
OsDD+D7dYlY2arD4gaPCws1g22F4S4wdIG9vuayMebEs9JgLyzMbGJgkwo0eVhsc
ANWgF+B0VULeTl/xVRYUzlMv9M870/QmMoVH73rrHWZpQ8dpsEpGs97tlbs46fXK
l313o99+jW1/tqlOndKN0myKjYQLpe2CDxcFv/EekUzMC0mf+RmJhu9oLctyD2RM
cKn+93YrE8sjpTPwv7clh9jLJgCsdKuCyanjROokgu8NmRKdeXhTcnt5guCh7iX8
yARC+Dfu2apQJ8clet5O7+Z1CI6HvHDZmLWRjDUEZEw4nMwhNNpdxbtan6s+pcsI
5N7ZqFLNMgzHRPtoYm2X/gaAreLUXfiHNx/8aOgaU1oB4726txHn4HqKkOHGOup0
N9R2LPDkG9QTOPirvC6GC9z3e4Br5YFt1QYlME750f0pRy72ATyUx31Cj9EVpXIY
P1iuNNYWF01eEDtaPAvJ+GZpyvd3O7/tmQp+75tEH22qzW+sb7h6yu3ralh5lTAS
/Us1vzCR4k+EZ1dnksZQu1lQnuMknAYJzBkOp+w0Djro85D5+UUllgmC8NcChfwK
JO9KxtyztEj8ngQ4kP6E4bvn7aa/MaA1OXp5r23PWSvLmSq/Fz5xLM2AneHYD76b
uGlMLZo9H2Lg6JsuhVQJfNlzzYM+1hNRD7DIgZcLSLwz5EnWyqAvMwuJ3VGps1zM
Q+nTrgplV5feZIjAknk0QXgdw8mbNbG0yqB2DM4Kq0ASZTWO1v6ZDdKdFjJB6wRI
SLqJ7vDG96uwFM5z60zPuAkH5I/CyBT0fTrGlABit3e9J0xnB2oHbeTbxBIxy9nZ
9/mLNdnJ0Kcpz5W0xTU2iuyy4HrDth6TRC+P/2FEiBrKgCGMt5RbAOlEuiQz+I5u
s+loS6SnmaiIidPqfxLBWIjzAcq+f8giWSOrBy3/y6KFSdRSiNhQ2piF1XHZ2xSL
b0Qnw5LWEa3M8R3K5wK3nQpr9jFZ3AXtVDn58FKgLVYi/15/T7H8OOWydMOgLutu
GTSIlciiPwwNltevSEOcdtYil8Bgcgg9WeQtAIFUNNI0PTGTmS27oW22ANeoT6pg
pUim8hU766b+ABE0yrMD7ayZTChVt2wO0g4+0u8rKFGiOQ76/OY8zK1TWqZW4BJe
2uVyTKpJBjrx5YnVfsxAEgNn0GsGnpQ+lLhwpiIEPhnElpW/3mX846P/hcGIXh1Z
7EqKfXnjvAI8eapqWCTy5lSF89ieFlFHiwVGcffc996uC8/mJyUqfLtevSf45Jzr
nR7ul26T7Qhu1fLkmmG+9TDqTTpMYS0hy/MWcXTYD6P6r4NGziT6++hTpqus+x8s
ZHHnHn8KPqvuVAUGvLuoNzFjWGdlUqA9r0LUYjyBEZQx52ZM91hP1PHueK3ti9uc
COBvHoF1smbuLQdu13HNWHOV7FMQUKY+5ao0++UTT0/JLl/1pabhA7hUX6ImWYGS
p4Bn5YYmTlku8d0Hd9noNcUzGJT7dAPoRdH3qNP90c91rzyGUw9OfYm9Iy58907R
BopZtHRFbxZIY3yGzMkgRFxwgKeMKoa3yHVqwheLIqDTGEKL9PT3d8GwjFjYpvV4
vXdniDiLChbfecyI8XpvaZRQ96P9oaYAI78xBsg7+37xuNPNVVHanngc8daHPLqs
ErqbXiVvyADBjkvWZ7xNTokbJkE/DMS8hrXgIf367CfQM9933Ugg7rNGFViXGQBl
qTnOT18ezsPKsiOyPl1wARaW9BJARcnKJ3tHFfG5f/OlkQCqbUzfQaTOu7uAzn/L
VDJPMu9KHMIk84mlhq+Ni9AS5bjpmU7Mk8ckzu2EZIutTqdRm4P+HEuLNmWofkPa
5QgoKvCNpAk9gDgT1VUxyTSRj7Z8NpC2FPxiMdyTN0GDXk3qhDeRQF2xQloZCQmL
nQanLoW/lxepm5SBtBCpdHHE/v5SQFZDxEnZzRfayhddI5FX7rzKwwd9q25iEL8R
nRX0DT4xHlvXS8pX0V1aFf7REw7PVDESJaWOYEwHNKjlGMvm5sipd1IducDE38Xo
JT1P6hc6/7eWCAxgIRm4MrX4eUvEp3yguFzJ7TfJOnLhwZ+9//LNe6Xke4GhjNUw
f+uQYkv6QhcJvv7EolaD02ySkyNwz1PReellnMr6Tvtl7Ewom3U+v9dGPH+ksj9x
Ww7XZCNuiJcEE2llcQ95v/SEly5tl1Abj14wQIZ87U3ZdVIlFQ/gQrNpo0VjMhM8
+MfBqZxD7sig+sCtXmrltl159M6HybO/umf3STbI1RtVPCiQprqDr5EYDBFZd4bS
LrJFOTcbD9+srbnfEOQp2HrYkUPODtdJ+KwdtSi3b+S+xenffQaUUgxKIBow8hz7
4vWy9FQIp5a74xNkDSVY0xol1ETeUZ9BelDBX3qHmSoEJ4qNqwlvbk/clDBROS55
nDJI/YKoL+R29zNgDA30yYhkdldYvEpCMZRMgP3gVlssY+6Rjm3E8jFDhSVigh0Z
Ri41WB26eO4HqFAehoW/e0NpI/0YnFmHnLTgte05UgQfZB9soqGGv44RTKnGd6Hv
22KbEEbPfMesRx9dSJzCZ69KfodObBW0VxromHUus6ka8M2LMkEMcTX7HnOIK6wG
BbDCR9KhmG0Kgixk7gSdtupUJPa+gBjAyxEFXzFDH5RhQ7sav+TuNdJAV1gZNRW6
2sTpvzAlwGJL+vnoEOTmfBDmtSLYLfN74fOsEsK5Y2mZc702NrAwKkwsOs75oPHB
OGue2hJ5Fvkwn/XraDnt6pugYLbDZS8EbTTTTJ7zX3Gf2rdL6iB3uwhNa06plO3d
cFaqRwmp1NxUDMj3D5nnyQgZ92fgyW92u2OZW1BeJKJfyGeM3buXjGrJW3GfVjJL
M4LpPEtv9lqQDiJG0VRUoqcWrzbXCx7RFX6NAr5eBNo7FEcohp5Zo2KKDRVijVCD
M8dGPLPAtYxXKgowSxh8DGrn71579ZWIOngK4iKcW3wWS6ojSMoY/wIMZuVeKP2s
m0UDZkJsg26EjqJEGn2fpbBYzkWb8TE206b2rNnHShm1OMc7U2w5n2I0VxYt7ezw
v/zcUAzh9Z1131QmOEcPf5CxLNjhvc2pNPLKh35w7K4Vc9K/KtVQBMgBPyPm4SaH
Z3GkOeXjSYgJ4k0tplPX93Xj0YaniCTctFjmduIEDx+16we0AT2mgz9nTGbfQ9If
qwlOfmoj4e0V7JeEFpbJ/d6ecy6kfk7LifG41pGMYlFR6uOU1KEEXbmA96V/bbru
B/H44csAYw8eX+hx8eJk9x8QdgsLaG7ZArQ1k0Le1p1198a+9TR0XN8T+r4HztDV
xdmwhAg8U/rrQZ7mgW8sJ++yX0RqDWV13rxQ+0h6wKABASJZVQajwfKFhVFt2fnQ
lxCO14zjjijHbAwzQUY40xPhmDrUpHxUSTvS4zN+NhyBK70Ve1M1V20VKW5MB1EO
tI1plZuS1VK+HWlNSgeh22I0qH/GTRscs4K0TS2e4pPIcWsmGxJqYWFxYZzqpLl6
p3VaSoDxQDCJ7NLCUZBM69T2Y2NfIc14OrGaQ2/oYGIfkl1T0xp1+2rl/6JAVu9V
4aEX2gLFUAXHQwMaKxWMe7EcyE3hwgKMf8entYroIk5s40RjF7FCO13nK0WRbN/D
Al4CD7lXeRIgUAISB3yl8iNRomPb6UizIGS5fq+aAdT7EyclK3v9NbRHueFK4iji
OQMUcO5qj7qgKEqVa8kDF6Gkv+n91f4Vmhi/6sWTEhRImEbIn7obWB4MtlbJZ/uh
bJ/JRLW5iRVtHK/a5r7t7rhjDCgKHW0x32rvxC7Jrzsw3/QpA48C9+Bk32Rli0Lw
MGQT/v+IK/o1BixG718RGD8OXUITCAo6QydVTsSbCFwU54qcxpp/9vG17sJQpYfA
3jZSNwba5aS9VLDyFgcPb1fnu/FgYheKlsab39qEKmslvRmyQixoDJQc2j9VInkr
hO0ahFHAQ0kJL0TO6u2KYOQ89323IvGvpV2BcsU0UFo91bWTnmQHUjBuFJsLTzUV
H3JocaoyqTgKJAlkDt7GbUqUzKyx7xzdW/t3lQbqltXUejrhOjYFxZGCzpNk6iAP
6Y67V7aQL8DVij6Et02LJ/NT+mJYgYGxtrKa87sMLAg=
`pragma protect end_protected

`endif // `ifndef _VF_PIN_MSTR_SV_


