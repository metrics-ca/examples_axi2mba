//----------------------------------------------------------------------
/**
 * @file vf_mba_mon.sv
 * @brief Defines VF MBA monitor class.
 */
/*
 * Copyright (C) 2009-2016 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_MBA_MON_SV_
`define _VF_MBA_MON_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
EMP/z8KvBP+TzpHH3b06YbWJtdDPlQ+VIPM8Sdxek0QWZLNpuHuzpeu2esvx6zwM
2gwLjWLiS/V0Im1SjAl9+UxbDiopmivVIAOUIXfO8caxeriCtXCTy0gF9QNBol0Y
cSoO/gXHjnFDCUfQWOnrTZBI4wLcOhFmxcSJVaRHtsPvgEjnY8MRKNeL9eha665t
I/cdbQfAkI7PCMkizJmgn7FzF8IKgGY3O/emlEcDUdZ+MsZH0wEpg4kb6X0b4sXf
vWLIRU2LiewZNOe8u9QnDbcZjHIODfSSHdqUSRfkG6gjvJ9lyu1H3fNgaBmaJ/WB
E/SyZ6e1HA1vRzAzcqL/4Q==
`pragma protect data_block
Ja+Qe6OxY42FzRQmVZVT7yIOmDlzySgtyDyzfacdCjVevJ9ZTUxAuvrUMHloDILI
Mg8rCGcQHyEVj2Zyk4xNIBM02s24Kwlgi3H/OsTzcpUd+eIx+SsDbdVrw8HFO1b1
D7ZzEE1l9khfyKtQjB+9HGENDVtw2YlEyVH/6lm00y51PIxeK4XSYXY/Op59zTik
UTJ5qFHDShqOex7AfO79RJx48seQ1UcidPN+0py5wvzsUqorb7AFzGR6wEZY53As
TD/rqFpMEFTwTsLR3L98/ptRQGvdycF1CGxrjSdBHjrHBlTuINgmzBxS2Nw4fEHF
mwrYCkt/ezgr9p31gGfwgecWu2Z32bTYnL4CsHSSHTVY3Li/7lZJ1nEttq/+HgFD
Dsw4Llt40EmWv7TJXs/xXv2wX5IxmDKgSGfiGVmQeh8DfSrTrmtV/RFZT4YFEVQa
spGNaCmeJNwxmX27LvI0UKs9bqhbbywUls6aNQ3mq5+QC6ZEuKDRw9Md1+jpd2Qz
XnX8xZB09Ddvs0E6kVxZdfGbknbwqliSwzhH4FcoSN6lHT+fVPth2G050eurmGYw
LFhitXLQ7BSzQPZJCDpD5TZF/E4Zryqmet6mHMwQ3k4k5hSUW7YBInRSf0rpAnT7
2pPCHJJfkkVl1weSu8egQV0VaepVHUgWzLmBGY6heDy2tzWYywjdW9WdMrp+HHQd
OcOCF3Dr7ig8Acy94WNgGGgQ/7VvfXqK2F3IN4EB2Jp6CC1bz6MegzCdPwJj1RGL
h99gLHUIdDz/AEUSNItmVzSqdfmlL7dDfINzNREofNTazEVF8BbO99phvUoVvnPK
uKMB23EY+uWbVeOj8HipHOnrYTY8XnWKePnypUaQn1k+LbpEdVNtX2AkeCUjSEs3
lAdq7r9nhus63R3BdX+0JnrVsqpcJhYuNhQd/qTLHVXMeV6O5IEWcCsIsWUNT+D4
2hv5O4rw+v1LfjvioFicuSSPOq2CP3CXdrVGfhFzfSCiifpqSq4WCiBPVrItHuJt
VMOBPMMwxK+w8CXvA+ph3kyYMb1Cw4nOs9SGOHtOthnP5dB263NnB9ABuJyDII6l
EropoXJUuHu1QRL2TlgJ3R0tcgB9efenT4VMhT4xNBJIR1euneitb57mHxO910x6
+4Q+WcdwtEV7b1ptSq1+KXIEy/19i1BS0I+zJWvTUFxtaQ+yjopsibNaoKyXI6sN
GXhCGZGcoLvOl9wf1rtC37YOqu/tckyfb9UNWOX6pwrkN3Z6zzZ7nRBYPXoHksxD
S7524KBeTf98ss3T2PvKGHmGccoXuSMnS62w1oTnycH1RiWogY9XqYm6DBeW8Rni
BXA63Cs9tfYBm+ffnBTUPWDcOYmYtr8mPFHzVfoDua16t8WucpkBLX9oEMG/0i/z
dwfeVHEtZfQ6f8VTzIk/ddjARS1qhsmW6xI2Jg4M5MdP0oBVsABQWscLMYrOSbHR
w9Ra6iEaCyvo+vgHbJrAZD1U1sUt4fp8IBA6KsKYMKIRMsTtnnBsOJ23QwrjKX90
JqrMgukc7mD+XiJUy3h1CDmSSfIEZ+B9GYe4aKGHPfGJdg4I5VJNin+C0NQ9gcYv
eEUJ/XmE2OregPz5JWov7AnOvFPKT1QMrmRIG4/unhNwguGplZdbTZYpekeWaF3s
fFrbXCxrckvgucURyr/5ccV8nImUCJyKDt3UovR7xKon2b753TITu4PATaTdHFgw
8gfO4toTI5T7YnxA8TfdyR0nIk1Mz+yzn2RFm0k7E9S4fbYEGiN9qWiOGgYC2Z5u
dHxHmuo6dDoyGNyaVfbAhnLiPRYlADlmBfuBc4FvtM8A5/TYTpkNYifRAUa0/FaD
VpNkNprMvm9XUA9XunPkc6K2fo+hLLZaFTHZORB5mcFkP1WLN/unBUL9ljcjCO+C
+3JtHrsgfEKiskdCNnRRVjAlL/4NshWYSVGsmNm9ZJC9zMOwO8Mg+O6cBn1dCUtc
r5z8Su04G+JrrZnl8Xr14T7PfA5TkJ38M1z1NqYB/VAszTnkUfMW1sT3bpepPJM5
H1TbZoZyG2HBxOCFQko7nz7wpUMqJCsUBcYUAgz+dloxLcAkjlpwdQsfX9NXNhWz
fHs/NDXh5DxiBd0O6Q2sY4ttwG/DJdDO2tGIXN8RPTfFV5VmTZJFW+MxtSl8g4zU
mGXLal4rkdmzVt5drBlY4RY++H5pJn9yPP2OR+wDBNMFGEy4dGeSdlwM5Nu0IwBJ
PikaIKWj1QJfC4qPKiOZf0Io/xiN2dXQmMvhPBavNhg44oTczVR4evw0UC+v6MtG
O6RcBW/21enqLdIJzceiDupEE3V3CLU9hHcNb7VMD5q6Zgyg7q4reZv9o0vRc52E
gH1Af881AgssKeOW66p/zD442nuFBn0QSno/a39kVgSCrUvDXqZCGraiOa7aRoI8
M8Uf3VRK+AccCP46wta0I975NwtPrblEiE314jkKLenAeXQuBfnIoF507pp8xGrg
o6iCqX/U7SVxIvYAkygi6f+igJ+AZdsjCFiEuKAN8lmGuG8PdY3hEjI3YxfPsg4S
C12ds2RW030wAWqMvLt6W825gXvWhnmNYPs7u7PVk/F2m3zf4WBW2tl4odn/J0Q3
+N64ecTIZ6UXK17NVr4NV6smuH/njbtppX6ZNQArysOeCtQAMrrleFH/Ih7v6+GV
3uFHs8GlZCUJSGYi2GghiI3/ZH4NPXjCac3loq6EnTcqCEXNJp8LIobj4UU8VQ05
ReK4/YREIUWqG1oUR+6np4/lhe5zb8zY7VDjQEMpTYyzPrburOy4iOemC+P90vXT
ptun3yBJuSOFd5vAXEZqzaFcR34xa9DSG/Y1qgnuzO0/dpBIcyLjsgNu+gt2GtMX
7iAfIQwBMCW5n3qcUEe0K5Xrk7J+04O8q5SxW5reajsjWIvetl04V9llV9NjIkMo
JoNqgUz+bizyBeO0Y394GPuKMb+z6mmPzQytvz9Z+yh0tIad/joWTiVYUsJVCfb/
FTzht4L84VKQnJktGzvlcUICCt6EsTTMVmU0opHRckJmZ36PYUfHUKCncREYlrz+
OZY3XjZJVx2C+Ff2zrh7Viu/5etCnTVDFPlLlshbRf/+tqgpIG/wJfUsTjXOtk1Y
9V9R+vUsjHBC6fv1+yKykRp/jCKpqepUXlzJrTKnB57BsI5QpMZp27YA0SUMsLbm
nDJ4SSO312bpskxUFDnCkPc4xEB9HGSZ8PBXZC+7/06nolVzicNrAEp1A0ybcK8X
w7CwgmQjYN5LnbBc5/knzsjlWeKyDQI1bw7Ym+qcBKrvR7VnpouLQkOG4JfFlUES
xjVr7lW5f3eGjueCGToCUKsIUub6OIt4AWgqQ/IVGes+Ii2eC4WdZvp0em4kYNGQ
KVrsKfjJwPOEGgapeCKdnJPkz6W0AJa/Ki+4X4FdbMcY3k5Hw5pTYqEyQyc9WnbY
UB+H8OBYBtAxA+qkw+6lzAVc5X5ckp5NNZcnN6e7z0QGqpi8vMAeh/EMcQ/RiEzX
lr2/3lCCy3QjCV4E2ZVFhKC4Yn0RqngWbJ8SgaGXnCl8bytnluCxn6QlSVBUEBBb
QmPDoS3PvbmQVhFdjoK4iVQta/UWZB8YH9Xd5BXfCYf2bvKtCi+/uBqq0HwsNT5o
WKhth77mllxk7mofdk+D2jWN3AOYnsv7zahuy4UkeDHhAylkgTV6d9xoGcyU/+MR
O9l4+OY8VHnZLrLDl5eM6dCGjezKF9bTTFcU8DtFvV+QMZMXRT/RI2rMV7bwVAmC
OC+tP0M15LkMYxzuZjENempVu5FnZ1sD2v3KNVMSlEL4uT0wVaC5mVKsjmWaZ2PS
LiS2W/TX1ghJELCchoYb+fJM7ONQWK3lK2dD4lvhBlKkHVVPcfmikKBK66/ZXAs5
Urs0HEKWeUhRYRs2lJVzpVG1cI+Py5T0hQPcpXEaQRRbTu8nno5JeRKaqwxKP4uT
dxWCQ3rjXrjl9K5AL2F3a30RBMdWgGVZTS5dU07I1hdAXct0RDSLl6yttNwT3Ch7
GmTegGuyVrLVOJa429FpTRW/HTe3vwUVsikfqxQxUbTwIq28bl437v9a+spgB4Wd
KOkTscZ8gcukyTQyX3eFCYUDuVTKJt3fXgVa+xX5cA3m80FVitgOz2Zip9Ec8M/e
Ifwy8jDhERPay2fcaGE6aNn8gX4ZXPKO7GALcydFbwrXm3TsCK/JgER01c0ipJ/N
XvhqeHgpxDBsa+0m0afPMh6UHd1+PZCf0GxGLFu3RJ/j1tO5ne+wIeyizNCirG+v
WaZvoEUX3uoP/1xDNkY8MVISh4q5gD/8CxRLdr3AfgbdyNF47wnEYKJUDQDcI3js
tqdMLn9JhDg8beNPH2djGLq66Pz0+SOLSLD60ewijAG8Q+Wz/f6KYdvG7mkWCTPn
6IOSxjgSKrC1LND9xR9YAVwXMTl6R2ycPafoTdV0WW/tzzBy0tNppy2q8xX5ttcL
4TJpg8M/1LXnvXK3I+ksZZBlWyXAynvkr72mG1pZBGY8httRrk56jZnNHE7x5IWy
zM3ZV+UfUYYdldDUG0KbC0MAl9VMio9L5gsGP3Fgley9jnbzoDmwlMdv3aQ7mg9K
6HCdVrPpxcGOt5n69nJyY2UUA6CN2ZpQvOPqMFSm4dN48TqSlRcVZq18Wpt79X+Q
0nA8dUI4OYChuUfE/5+qJFPMEA2gb0sv3ZIkH6g1MnU/xJ6jUwuKLjNofif00sZC
eyfE8Pa742rln98OmDPU8cj7o04AeCAzLqYqt8Bs85OjXx+yKlF51Kd3YszZ9QOh
+FRSyM8GI74JtHsEqtcQsDQm0L5z3DPZCBceOtDjrbRcFL+ScJ4s6q8R4BUMvG1y
lNy6hADeEluEMPB4uEZwBSEI8fSBljc+oVZ97u8JMJO6pA9QajOz3ZkDZYzd1RqD
eKyYcwwpuaoQXWgmlg9pblnRbdQ1HGnBY64x4i6ib/Mgo/85wPWY05vlvtPym+g0
rKweKqsenfag9m76ObxKFlcv0ST6kYbzLmds2ROK8b6vzM5h4fAufz/ZjpzXxs4h
eoNpAg50RWjWWvIEd/vHjvQPWBIWn1/hnHQKTX6JkIPwAJPB1EZ3lfVJXBbxh2TJ
BVsdvI4jqQa/jPfXnUoujTkv+Wr72i/HE/XvaBniBGP4paztsSl15jYK7tO0Ni49
Y+cEo9NiZX6PxO8PBvdN3Bi17ykDvUbPe4V9QZxRgvMyyWgdkzCwl6nZbiGf/G9j
w9onL4A+1epbfqh5cYeVWTIpGjy6jG6Wy4dq76c3ET091+kizLGxH753SI6XtxyB
EiGF9hQTXjBdIjxXv9zk0S5yboucQPNsi/hWkkJ7mIm7NwqTwWN2vh6CDlbaR4I4
8SqBA2S/NCtniv9/c+NOM7wPCjMmCJHzqsZFqKz2H9O+NINOOO16jwOGEhzKnYQj
uj9VyIpnq3Zxt0Ir7WGO72Bm9N9tBxQ3SpbEFKH10WtsE7hsi8KbVujDE9yVYYjE
565ZBU/p/jp/TJeQTdkxx7RUG4JqjIRmvNeUuI4uOgBLwizbrDVjO6ZueMboWlBn
toLxT4RcOb0Cf0ibiz5sL4fs6UGNQj6Lbf9Al18SSsLJzJBck3hrl4YhCqDoWHbk
KoJ7IMoaqY4Apl3U+xoxpyRsvC0TCWSH7FWqre14MejoQYNfq8U6jhD0wQFQHquO
nm3f6+9AWSGD9qXRFf3YePDBfMM2LSiRyT7CTn4JB1hqOckJXiD1uHS56SAhZPIL
+AYpRKCWzcZcTcKXIx9TP7Gnx/+koOa6BLZgdA50tGNPrkCCTWQsoppEw2hPzXrL
X7LtaSY19Us6QnLZ2LezigIzTGCys/MSdQNvlzRAzeit6NzjeAW7s3FMeE8BX2Bb
SEAUEe7JYIuSjQyCoNIpzY8DNzbMrhU3oj5PqnX8qKmr8WdLf6AzCClrP76pAAml
Qbg82dXUm1YXzm5wrRI3K8bvXEXh0dEzKxrWM9LzH4rTuov8IR4GRSfHNs8YeZsC
Fn6jvkknUnwGQz67qcowGvf+q5PJKP5/atXbtCXHzXyDahdCi9EbV4b76NGOQkIG
HlqAlNbF7KWjw5bgborGVbNpLnQ9QHWJSxBCTMKs8cQ0b1BFXeX+540GUJuwY+8m
3/N73vQdDwbo7gxFJSQFjL/8Ej1Ru8JiHQbEYYwmvBRiL3znNDRmFFAQMPwEy7Ji
BbbgqlwQJr+jK1ure9pnZF5M7kG6Y2wI+ywCmpN/Xktl3jGVHJQWlJcJ7EG4v2uY
B3jDDGsz279PzwSJXsiYWd4h/Ar++j3MTJgJ8R1qaq33AxgzmRGdTj10GfYMGQ8p
5gzMGLeUgT0IzjwDMf8BrSQwkvUV480aQpclKwc0tTB9AAw3hAxizeqpSDGXNla9
psY3z+Wfn0LNp/W7LRHc6iLea7vvyZLNUEi7oN9dE+DZdt/aFSXEw9img0ZkJ0Vn
lbHbekDWgmHHEx2XaRKKnEx71RXvEeFpWDOq0aI9xvVSMFDFTo3JpMkraz3XO3WR
zgd1OeBKMn7v3RVNPUiEYxMqVxy/9fWjSfgeOxSWrgfkebuBgqsaAS6kOtP96gml
9eXTZ5FgxI6zsmG3RNhA4oVTt3k4B3feKP/jwk5lMKLMYtdINzHR59MyetpAxAwt
auH4n10l60Vbh3xk2y0G5ahxF/hNc/ikgCcJxndn8ASnLsDcpJJExVl1JNin9jmc
wCwPcPRws1KP9HlqYrWpPhGpylqh3c7/giK1u//4QyjAiK2J5wAc1k+2NduOqoa3
Lh2hQTYQSzIJj6b1ox4LpS6s3xDESRPGi69b6bellJrxeChrTI0OcEEqr46Inh8N
OgffhbPtElxZBZrLIkEi+uVZLMIhP9VU7L3HR31FLFyJJj1C01eG0Tydtj8iWfWj
kkYZU9eHxR/0gyISu9r/bLT213CAxapBcsqgl0vKnigQ143tq1fmz2RX28Fu0KbJ
+1V3deUIztuXLtWX+22F0GCXMglxOH23CUJnXF/CHdqPfuTQY+nyzPmMV63aCAgm
bbp/Hco9oOtm0xyNLVO0jOd/oM89zZbzGfYJxZoZHvJgwUo9mx8RXAQ+uKY4kjqP
FyDI6+m838VcOB+g+v1lmndzh8swEA1oUtLPnZHeqw3f61ydjR973lenergsujWI
2iixpfNsCrG80a7mpKnHLUzEWJrHfUFV68Oyv8B/rS90oVxh1nGlwfv0ZM8WrDp/
nBss4YII7EIf2RnpYp50DD9I2Kejo7fgsSnhwYpl+16mFrQlRHLFXFP0MaQWx7B9
FnPv6bDCBfGmdBEKIRgR5slEiNlLjpMH3idQzg7Zzfu+mwnBvYBmhUQXRMjcVrT6
oGwn7tsHX8nWcpgHPNAM4EYEYSvUSXrQT+S+j1ijw9Xd4IDimd7/B9wa6zK7Rglc
7iYQRvE2U46leLVCRB/g+RLJPnJ3V7kTxXqqnPkThzFhhs7ml+5UW4GPJVEvptcq
bXF3SIgIC66ZyS5vhkhcsxW10Get2Zg/0oQeREqYnMEpcerdPzkB4bcbibu9pgp0
Dk5mfSkFtFo9yD+ZqkESoAQL2TNVj3XtAwaR8yaTZbrZARrKA4kfacfmhFLiwwnZ
UBK9dYQZPImCDsWseyfemVZuU55sNHBYWiScap4MAt0ao/UfIX4ZhG8+RPXSLJEG
jBvAWyHaFFO2jgcsQeOuFmSS2WgnjGq+lUmrrYPGey9xOcr3inf/q/wnvnj/OCpg
BVnfTuHvhdUY/6MVrFmYNrg6d3agCLmnxVvcVB9Ei7WpfR7pTdBU9c3DWcrl0aDJ
FmuNrJIG1qsT9CCXnyH8vV0sKezFGyUXBCAI3Jppmdq9o6wIkZ6J5UvvQ8aNnaew
kQd/bU0uZGKeKHPYGzQsk5MlgE/dwnOpcZt/5O8m3qNGrwkgc89eRstaeVEYYmgI
ZQdeytNLhMSZV9c4bb7tWxrQ4WnG7gdESIM33T/63sf4Dn9mrz8lcCMRm2Vwky24
9zrUMG/6Z4+GOUeDzfLm1ScgD5T2/CwfJ7aoJM1fda9zR93tcpQ+zB788Gjwc/Tg
+d+3Vv3sBZBYH1bKVb7WT75/ykaLRDkfdVtjIl+r5bKAMZP0XmKMSW/jH372D9Ep
vd5Q2w9akCl2cEjM/NGaK4dhEPRVhsNd6riVhvNV3Ghb9e/9mx6eNt4dT4vt1zXf
wAoXRSfIx9p20magEg9TjfUAHowNQgVZeFLLRhcq9N0PpCcuiMqtZE2a3KYp5UMs
jZJzPnN7ZeXlBFH1H7UQq2APXorzU6YyOY+qdjkfbo9R3Bn3Cu2Ga/Mdaz8/fk5K
gNrId818QQVfGxfiqJzaFiTN4aASBC/dOUP0JVe7PWF4QCDl8XMj7JVo0IEBfcqE
ZulUr0UKvCyiXkDDnYdSe1nWBpr+xdRkRvtBrJgFf8Jbb0CjpiRfFgDonnnYq8SD
RQnrvsIroA1eEaUwQ4W+V9rjBfvFofhNQ3X65SA9r2votM7YSGvXvVFeuMBqpkct
2wMSRRDUthUU1MjV39wSdrguL9ptr/fMByC/UK/atV8CLgvx7c5US2rDYmS8fmzb
D9hjPKWfOidorMVFoUhHOxUeknUBsxdkNSBjgEhrSFOARQl0spFM1o8iHL2qJlq6
yKHLctfXtGWZWewNCV8BzH7XTO+9Tcm7eMjWHvvPo2MgN5aLJZ7Y5K2nX/ZtBji+
tA4kcRck0tUYGUxNWGTbndaT8fFFpQoPAqV9Fy3/Bpvnutu38uZWRKO26Resor22
ABxc6KRj0v+ckF6vIgPumd4BAuMepwEZ898VnFXNH2lBXZuJNW2unI8/4n9rHMIF
LubQ44gMq3gclM1lqguIAnUg13B2eoFCLfOx+WSLdfHrRIzW3KukA/2fBb/IFQFd
5zluq6u2icKsHZrRarNzCHQN3Fm91kA5bxVNwZ5/ZblmqIJm0egRAlSWVejFUY6R
b1NO1nRGTUO37DmwM4wjHMTPjS9qMcuIA4lVOIftiq56GBfhZTPCH+NikW5Z118R
nABdI4CD5CzJNDzbLgFqKyqJgXD49JhmyHtRP/2o/PHaF4F7aopzHubKBegdGvdq
rA6HFH0iRnP0IUBBVMFgYAVdya/qT0Cd+5dUI21qIq1DP261RCd5h357GcMZMYcT
xHvg/fR94vRJdMwuNzjdd0PJgvBAnwa/LNXObcykmcq5IKTN3O8H8a+YejTnl8CN
qab+2otWz7/5k9pHOGqmOKJoHVCXh0pUqyQ3mMAw94Od+5Xd67u6y0A96qQlG1Yk
D4s16/wQxMOaMEC9bxG4HzhjaeEYXB8GFeqKCrhJpe5dNvSIwmWRbq0C/NqUuPsl
M7gpT68kWH72HK+x/Ry7mxZQH9ZjLMiOuV6nh1rHzIKne41DSvuXHCVcYpbvgC8Q
HbRpplmkqhacUvUfClEK/tforjlmOK72tmVPkGnnYhvWyb8Md26V6ZoTCDqsdkWO
hNQ2hrX9OD1FeQoNExFyrBPiTzkuVQVimI7+GxTJGX7a5wGTP3LBKJzSi9UizUGt
wHjSH8A77rAjubaj9xUh+Yf86vwc4WXzaPTOHYLhqmy88dMcClXZDc1m8UAHtiZK
34YbtdCS+I5F+563H6qUSfPudg2yGIYA6n5X4jpFw141JQzNVpgl+mxeNsXZ/oCv
s8uhc3jaYHzbvMnF8UUnvOWB34Y9hvWJiMcr5IPCKNrVNbop3XKt7xJnTuIKXEfF
6KNqOiZB0M4mGN7h4nupEb/w9WMIvZBbxTFMGFC4OLsF/coUNo6OEAaP4IBNsAep
j6KDz6smx0aOQwx5miP0JwciVYCbQIKFUMoHXR/gfU6eQEzboTm1VsKRhXUDLFlr
4eSxaJVD/pqmkAbh6xerOl44GN/Bic71Z7PyyrXCKIAIyyAXUNmdRaOTAWXkOlI6
sLsXktlM3GIk/zOd/HGLmHP5wCiVVpDTt3oa0WEuZZ3/9JMO1mMkU9GNqGY6gKJ7
7eXieiOGqieO/MEZfkTQ/iavzC2YZ3MCy1L3Au95Kr4vZjfTJD23naQL679i+GqR
LJZ9DnnkPB1uDr9hTEtvexZHxiXTDcHjECvg+B6P8myHWLjiRn8fuGKENsUgEuQD
NFk5aYLGZM489uS6i9rAsygB93iZDkITAEoBqT7RdeJb2gxjCrtRYY1OP8+PPIJM
UAoTEXADgMR11QkYmcovXYMHstqBBGx9nFZ9B1WjgSb3t9m49uM3IR3CnkczGweB
SkaXz+zprhxNEqHPdD8Gc9PUXSRtBf/9j4sBSmXo+puqFo3Vr3a6khTkdU2pcocT
B3V5/du+ZEA9rMJHzEnAUzAfHcNFtZdY9lvdktaGW+sspFhBtwzBV8ooBSRv7+zQ
cysavFvl/vrn+BHKdE/np0c8bEZQShpgFrE0j6xV4qwfOICfrmhhnUa0b73Wq3Sa
FaeLA9t3LgDC/0tqvYzWeLD3kFi5NIe2KT/rqTHwSPhxDK9bFhQ5iXeD5Yfb6qhN
bQ79Ll2KlVTwncsefkXnh6sXeb7A+mhiA4DY9KThxH/SMTQjtH4PPgxYnQNuvEx1
IxBz3wOgmLx5VC00qqHBmmcU0V8h4wK47ssi2sl1kacPWwa4QVunxYy79UaBE2LO
n3cml469rwY5ujOba/XeDHYZiqy4iXiNpBXfRLUs0GAD8LilfNpeTYOrr9wdqF7f
MPtss5NISKOhtuGxJxkZdiqEQTsFOqQNJIuMouMwnA/OOFTMwiF2kp7wAPnsQ/GQ
5Q6tJbSF8Ccoqg+JiUoBUuZH4e4tHfub6jsQ+iZEQZuMswllCEbwhg3MQ+5Krcml
`pragma protect end_protected

`endif // `ifndef _VF_MBA_MON_SV_


