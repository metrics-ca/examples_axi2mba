//----------------------------------------------------------------------
/**
 * @file vf_axi_xact.sv
 * @brief Defines VF AXI transaction class.
 */
/*
 * Copyright (C) 2007-2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_XACT_SV_
`define _VF_AXI_XACT_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
rZc1OTlZgJc1PgPUCuYhad5JyZGqzhWQfNke3Kft5qjxxDzenr0hjrpeuSj862UZ
piM3ZABvprw69rBlPb1yfbOTVJblVxk+6P7R5Kb9kCIuRqMRcGf/CrL2jXwKRzcb
lPbRGdjidyEbHixBwV9slgfnzK4bU2jjgyVOH1tYcIOxLnGYZ/Ml/tEwuNGjl60e
+CV6KZH5K0CUqGkcdHDw56M5gkoAplXLbVNr1ecGn8cW9tGhbe71SuVB07v0gqme
ejiJSMa98uTW9LMdzRkk5d34aEHNEeroPYrm9BTWHv5bMULhqyVOKbPoBjvYbH4y
w5D0dJw88ZHq3lZ4obaLDQ==
`pragma protect data_block
A8Y/g8bhYBzJZ2gHUQMA+buUeFM7/hHoNIEkooew4d7P+O2xCVQABLGVqiCzLBep
Jw1kw43SznN1JEAjPYFdlGI2bpgGgro483+ldX0aSc+0PsMjrPcr5H88tLYP/NdF
21oVSoNPIhrDldgzt0LyA3ESsiJt7zq9Lpxkqzw5GfLmo0cgLcweaSji+xRrBHxv
VdW/XQD0zl5Y8yqGyb7B+A4T2Z5VkG4sg0HhSfq8XZ63JcKjhYgv23/HGsPT99JW
2vLD83vfhrkhO6QI3e++wN1c8AHitJoqbbkiQWmqRYt2Rut7F/Gt2FTHHJVlZ0/9
HGxzwzcGbat8AHAaHZAGfsbnB22DV1lLVrn8JCk0FzR6XrwxQvbvT/t0EB+Ht3hT
vp7rRoG1kgDmtBGAH4nqCdbi0Fxhj4zJ8+o0YkQVyF19PTiZEjprVHbpcbwdYfNc
AValHbF02fimexyznkl5bYTxKOp2a9NmXrD7UAc9wkGUZiX9RCd9PJZxNoWA3mI/
sp4coRq+jdieZilhs0QwsBQhcgzOFnBcaJrfFUzccJAlId/Y1GWwfKes7mRN7PP2
yafA6xRdgXM/M/n9uO/N/mgomPUtgzkCCKrUPY04bIpsvnb7ztLlleZSPmTLp35H
FE7goht+XhOSxwgW8+rcefRd5g/Jgroy8/G7n5PFhlDZTRelHdkcihnrXp+EY8Fo
dJ5tjV5FJ88e1g4uqS8TNtDOsPa4CmM6jCDnwuUN0tTZRhsBsHl8szfMwYcsV2pV
ddaLOmToQQ4dSlXnQePQyy+uC58+uCo78EPA3E2BdaFFCNRaGUti0ZEkoZUxhsNk
r064ABruHSImW7kZ0YzS8k22/0eyaJs9DtkHl9qZxAsfy1+pCu32yIJCy4aR8cP3
ItJprSjzqam1c24L3KakjmeGcawuJypFkjrnerZA3l832SD/GEpw0gN82FjH7KtW
OkRzK3JXy2AZ3vtmWTkdhP3cVwFS+dV3vSIm072Cpe8qpU6ploWZuqyNx7f1C6mn
Ulhpovh3hapINFs6rXhz2H4nWjRiYx0wMCkhY1PcoH/EhvhxoqTfEBidUsvTUKgM
YAPO1dn0sVuGqZ39Z8oXj8B6t+n87cEBYrjOu5w2udlwImXTTg2+4GlLnsr6qCI5
fsRg2648rt7gZJK15EPGuQA5sADEwDlU8maOYrBRZrPh0cNgzUR+ULt46Xj0PsT8
KiehxzS1SwJgl5tQB5eRncTtk35L0Tex0J/S1bL3KSMp7oecE8Ub6IyV0aw9E4u0
e8yjO0Un1K7TEerw3fuq+StxrsoB1asxMxpnicCNLAkS+GdG0yZKU6Ozwewj2qwp
QuxLfQU+KzudhQz8oYezAxlbvNRhHgjL4Z2OQzsBiWNvgw9auyrav2028pDRm5t7
SQx4/K4lQdesD+E5sdb/xPlAwiEkAjH5VnHbOJZbGUhPTBKy1YwrnKYKsCzcwC8P
6Z5FOZHX8yJURl7eoucMxgSHAfg8sp4op09n0S9d4EZVM2rCBUwywjCjZA9U9Ogs
Ns2rH4+BhDgV3RuXFZk/ZWP4HauZZIPfGvUnln/FV8AnX2moxTwYiTuJrmOmttEq
nZuFHWfzFXTX9eO4cRFXL6P6CtljzYhgYF+ZYHsiEHEQYCzQaUCJ7TTTRFtgo64T
EAac+1KCNFZ34QpdCJ612Hqyh7XLKZXEtpiNvvN+H9+iFwWFj1nzx9WpL+B7fzqe
S33d0pt3esod62gCb+xyJYU3jYw0JyMKjahJ07tDfemSiYGRH337DxQ8YrrVNVfu
mmq1t+bQUWn61LXrRW1Yk11fEl3N0BmXSGp7rDGrZQWiDozEzaS9FoYSCmLsskl7
PDxF3M7vUvU4Q+Z7hdP4oGTQ2HgGLyb9Ow45jGcFZX9MpxQNdsp9KGWizHxb34vn
r6140Ch8yuxYxaB/d11uUCRMjes1dIXza5nma09y+B0S7zaXBaj99mcw/KProViF
NE8WIx5QRyKRhNI9VrB6CQnCTdxGOK5WDPuTwsRAjKzn8dmzcDTxVF9FgAsfHBTQ
WmLwFc1+nAuXVrB0T8J/z4I6NzWLVuR61a3BJJiSbBAPd9ntmUogu0YNGWB8IrsS
MsN/ycJR9Ou14AUmnfl52QOMjeC8wNosOWM8VaqH2vRbQYbXkEE0fd8EpTm5S59e
jeQvYKyfmK/7rzEiGvXdOKsmIJhCo5ZFaeAr+O5CNOB2DSGRhI7sstXTCAodUgJX
zW5t55ehb8NgJvXsz6iMxG0E5bKQmK4PmPWTh7i4xt07l57UgfjjS4DcuzFM+wn6
VlYuAJcq9tc+OX/YM1i9z9iy9aLOFR2VBn2Y3AyHDRBB1rxdePBe1TZx2MlOyBOs
O1P+NveepbhzggStb6L4EtMeGgC1MhI+vU30m7k/11uqTd4OCOZj6Nxdo62fvfXx
xR5hOlVoCp2ZggKJvCpzEB7wh62nB1r7pXnZAWxVlbuZUyRccDhL5gbNCrRkBLQC
kdyEFqtYlN4sTFhHSyjsQAKQik3zN+gBsjpGzbtB7+qZzrc22O6jVXGvRu6dMZ6I
Ju0UW3rMhYPQovCPd/WBBk/hrW/7lfS+hmG6VH8HcU773oI5JyGy1d88iXXCpTzj
zl/Lyy+WR4TzwsOG8QDQwDt5V1/DY1xBECmytEWPhZ5e/ygOdN8pO2KIEirFfgNi
CKGPFvnkCyvrLU9aqPvmvauTG2yUR42m8LiSMe1LlkGZufgMaLWtFQHnu7It8mP1
HPZFv7FXV/n4HzUsqu7VkbQuWAB4M6K19BVi+qz4aDMW59EouuUHayvJ0cBewZ38
5yyQiPOEb1d1iIcFsX9VwHymX/X33jc+gBTPadPQUk3XyXIeLutF8vZJTT1Gjuin
e0JZ1xpPyKdrQC8HacyxkNgVCPljYnHVfekUvFngqQbXAgIljPHu+UJ7TpPGZ61z
u9Io8dLJFF2j+OWrM7M0TZfZLrePbQDBCMUlHBHAXGq45TQJPgCga3wyp/tbm16t
DMwAoIRzON/u+ElLFwSp4xM1UyGK7G3rFZdScSor4672hvmuzrJsRKDtiME0+kUo
0FAJbrbyhXBMcD+a42z36MspV8EJAWVUjCYIorGv2iWE+8VE5qgSFSD1X65OBs7H
GgeobYeniAI1QKuz4oMcGQmqu0PttyMtpRmf15XQTVG3d4ARCuHlBLOkbfYktvgr
QHIbiWcoyig8ufEyjFyCzJK0uctt5+rByVCnw7KKHcs1GhXvfw2Pgb6i/uXVzAam
srFVHlw3CFagkX7ax/lcGjIjIyGnqfFx8kqDw6Rw9JCtxOunvNDUs9pxydrjHT9G
cynkSsrEYjopmuBbH7C5fdTy5u7CmEJ3Y5/pHiuDueBa7dhvjl50fIQ2c5D877ON
p5D780R1p+677rXsZ5sVbfJD8ShcmxPsqBoaTPr7g+9KQuC3eMHheq0zIVUPa1qO
YPdy81CPkY9b0CFYSoVF3XqcCcsm+CpKMXWq3gR+FjT+X6TnsIhqDoebH4N9zFvb
Y9qGEXzF3gpkzEamCqU7ZUdTP2u2dV9Xwqivxk4Y6zGmso5SB6SfwCg6PeR9Yc7Q
hhsrzvlULejcQ1VipdW0HvTdD4TR8/Gsb08NPrGPxdM6cYsMVHHohzumCvqzY4zY
QMZ7BRxRHLr1e1loS85gcFTLE7HtdMNTH1yG+oe+DSivozrrgnm+KoiTpxfjG2ap
7kqVVwDtjrE/DbSgWMK0elHXakbH4Fc1IEloJXNA9xH9m1rZk5djSjiNxtIx3NQG
JSPJrBrce59WoO91nHZ5IV1C7WhTS9qLUI8w+hW0wTa8ThXHtwbiXxuWxStMyUYt
G8xZRs9IuHkjpgvC/9CNRLEu4rtp00+jqmpFqlqwkBiDU8+Q/eb6+UYsm1xciyko
RQxJgxyPA16IXEWLY+OpPurfDfpUkDL9juz0Ca/JMBvdjGR0KFegJiY/yJ8OKGsx
4UBymRony8xcJOMXLHVhn5Socba5u3NbYrmds2gWseHrLtilEWjHgznpdOAR5tKh
LdYdoJIcDjiqzrKVzsNMBnv2Cuf2GLuhpbszXPk0LCo/35oPy+caw6pC9hWTPl5T
EOCwjZd8MLNibLHAfMEI9xjtLRQBnkzLYIlJJu1rqIfakNYSj5e3PcD7oGymq1IL
+LN8Fp3WupvslXHVgx8kEjt1+3yYluYgCGqJUbTYz6ItlAqHvyc2N9lxAfDo+kjW
YILQf7CEzNwJI3v7wOLKvFaQWEunrkRZlAWAi5G539NGAjBjHVSjvZnklQU/ZXMw
KdvwM8lU4rDDNYVFXDhCCC1iusgVCrOSF+kmfLLI3mXPoFA7BYSP3uKaC0bRZOC3
gNWnF4pkF8+wxwCRNRbAfiRuNg6Lj4YssCwrbkKRUcoBpkz11/ASt+InVX9BXWSL
o4+2a/MBB2787PXc9QQlvNGk8xLttcOVPPb+kM72xAkNUuKgblYt7FFTZlq/7JJx
jT+iRGomeeYeqBOQRDToRV3nxt7tQVRT/IV06MXl2AHM4wDJE5McZXKCzUOpE6A8
oTu7S29uvqbRaqn03FNjDqwIqbGJ9+1BOwcH+fwAJ54AhT+lgYvOqfdxgXXlCzZm
HFKz7a+ZUyzfJ3OIoMI60Q1xIV/jBupzzKsNhdE9a5mEq1FwKMBd94D0+m+rCzy0
Ju1aIuj5sPv77d1TbPNAPYSJFvHdlxWcflG7XZM/GElXHcSIXJwfIPZ1vpkPHg1j
u6v+JDNbBbGfI3nSwNT4j3kHVDFFiIlek8TnN6gVxA5zJD2nyiTLYoSLoVEY+/gu
gMuZ6P80RN0a3FXONwDwF6GBEZt+oCGwrmSDd92w0eWosBToZpb58emvU0IAxnCz
7ySxWwa+pFRN0lTpfRwsX8b7E8VrlPyqXfD00HT/rycUomorSe/1wAhHcsETBheP
fw0Yr6hxMJ/IFNa937sI4Yab8cKOjGHrvz8t4ur/c0hqGAQ1K9xex5cXtT6jq5hZ
NG7Fsb464GtvflMzAKMjzuSSJdX3de1Bmw+J3FG55gCJCmpw0VVybOK/PECeuIXP
HyIfrYrYfs5VcCOlLJ1di4mea+uNNV4WFQeZncrRCtYGGDvX9od7rDtpXRAebYl8
5JMgkLXWB31fJBHbq1zARvRi1I/Tyw5hV+tQbTSzUfU9i0c0PVGiLQg0JEKiBYhO
VbaAlvJJs4YmXMO6ll+EhGd1jtKV/wkdY/RBvR3k0ECUrrmQYswMVID5i6WtVd5s
7iAUVLvlNAsB+Wp9G7x9YogVR1qSXNQV5IMILoRi2QQBa16klorv/qm2gxnvyIsk
UMxF6gFpyBMIO7W+VOExGL0ZlXLLtJoZIF4jZKVt4NxEFl7XE6L4QdLQq1iXib/z
bjFGgGLBT9cqmFrJDEIg/lax1CZszgLzY2GcJxhIE4T94+xzBxNFT/OicYTgUrWW
d1lWh7IRjFDPR0lg523Et9mfWXhMaURrsHvKMAGSCt8MN+YPA4ELssulTXHWw1mP
FOl9ThuRab3ZgTEk00kQTE9tji+VtwYbjq8iLDfpwB3VDla+vDPZxH5n+bwB2iUp
tWY1VH8yQjO1x6GUbDUNHqKBpQ4OxnehpDjfXNjwu4qa14zEC5tnFcB1zvmqCcDG
t/bRBVjzs8JIb9BIxHFS6WyrVxji/0IL9TYl2m7h9y1M8V3egcdCYZEsUx6WDUu/
iB4gFbH0SnH930LAQK7fsC5KeJM0D8tZQq+duJFxie4L4xfqgnQP7o6TQeO5jqVm
HNZwKTMdgiYDi4h0VwhAst7xDT8RJ4yWITRNjYKjWBGXcbNf1obqRYwPEWm46bAf
5ezgvlxb0nbtsfdJOXNPqB+q72jUQzjnrzMk0Gg84joKT7NQmHpc2PQifvwYWk5h
lbivbf3mjLaX4MV/jwAxNYsQ1M2VyD8Hv1yB/c1TgYmip3K3xBcN7MWmZAWLMqs/
R0f8lW/B30CPOSqSnC6MPentWdcWyIVEASLCDrWQQnYy1q0dst88QbfQZigJY2CR
wuQoDMAf+FNTNRMiNRUJA5gTRfBfW6RM7DQzgJfVQ+IPrRn9lXPTMR68DC4XKYV8
DXJXT3sL+mhEm3yI6xXZWcD1qGhdxZfe6qZF+fXv5DtPUXxM4ZZmwQdQCQXWXq/H
4LlxxiFrVyj8QN+MF6IcrpTMu8aK/7z059L9+phwppL1trioi9+OmsnSDaSzJOib
EKTG+R029aw73Oc2BdiZXYRbTphJ1orUt0tnitFqTsmbvVSRMuQ3DijF+JXprTf9
CtmU6x3knYcYdT17Z9UC1CraUHV0Eq9ErHRQfKODyhxIpZcr3inEIY3NI7f3JQC2
lJ8AOLWvk6ccKeb+NT8jJZb2/kdqkGczPYvIkVVvBA29eZYbRf/aJUYWAn4Qqtvo
oQd79k0LdmiU5b+2U/jMh5+SMuQ6suW/XyqZLminuymBZHCLANbrflEybKbtND/J
Lz6WEbFcdwweB5t/oPcFNJKd+kC9ctzFXvdKS814RyS9J+I+24DBgExQeC9GROWR
sS+10E1rUOvPfiUNVZKkzCrl/xoBC6BO342kxC4geRzDqzksrRGXa7UgAlQPzv1Y
3ZFU50/YfLqyEHMvXZepeRTQeNNjHiOsH2J0+Ix0djr4NiuGx+KN1g4widljI+Zy
7MxrvoY3OU0atjCDnJF2OKAMrXUD+I/FgwGaOIpEz7JB3BT/Mj96XenVzFxXwRY5
lDYRBCXsTuFVzTLjLtR2hnbj2ITO/Ry1NoBeZm9u4Aspjiz0oJQ2RIBvKoZYL2Hh
HissMfdrE+IE+/ZBRn91lUrZc+XZ661J1uaFA1qiGeaM0fmU6FXkHNP0svEUf+wU
JAPJfGqow5392cjSuSJlop71DXiAPCSiOt3g1SEVjV85oeWR+2Y6vUCecp0EfXqp
RlZKg3laD41Dk65kfzsKMDVB7Cyq3ttg3qBHlNBWB8prvaLbSQERwQFys/AoZr+r
z9NkohWPMhV+QbwMT4fhKEAOhljMxqKwOkUwAFyrt5a1UTNkJqKTcw4b3+1axJ+c
lsaHE/qVbGy//ItF1zyjxauD6vNzcTVuR4ZNgACNfUtwMadZfdN/apFykGJPMtIX
YSOh7Sy/tr2twPX1Vrg348nG0Li3h9sjA+hQAIZ+KfMITVYuP4J12d5w4YAQF1yh
BYG4Q3YFHcqFN11g8hG8lG/ahkDwgUnewt9yNRvB6HVUCb3jIFHB9tRl0qFSckoN
GSEF5BICdIB3dvz4tzJd/UDy3fwf3H15uCz5LjnfGzPWknZNqfV8mAX2YBHa6VBb
zidCmSFBv1QV8PSx2/VI6LJquyT7rj+kDhLIorAfej0U1lwdZAhGSxR4L5lr1imh
FbKj9H4bnMngYsAxf38scCiVk7pxktlMfVSpevGjI69wuUCnTLIcXbAwM6bMCsi6
KHhIJRAkSXRNo7CdmNyMghpE5aRluUREufUH5iZDCwakPpmMQ1J+mkRYlCYXuXkF
OI3tlwTILROBlKGT3MYhJTAmkYMhaeUai2aYehq5x8nLdbbFqYTSaFbFLTWL0zac
m6mVg1x7GrjfzsadXptXy7++sLnkmQF26l1LMl07h4/lodvC0OlUbj6GVCVknydZ
IqbKEzxgqcGpxgktMzPDkbjMuhIY075Iy/hoV7JH3U2lkSyRklBfI3MVCCWsetoP
Ls1OK425qRzvgy8Bh9XF3ci9A/2AfRA+5BRTEZoD14JctyNmtTfnYcE/5+4f9jt7
bde8zq9t2oJM0rp5K5MAbc620tpt3gmTow0C8grXcFZ8JnW5MVfqE8x1IcWhJYyH
wzof3OFvJttwy5iht6H5xLeu5eTOYAzFJNmSzTSoh6hK43ThL80W86tcAW6VapP9
RvZMwee8wdbHWaoM4JlUHYVD/i6tC4Pqq0u7B8WNHO0bjRytP7w8mhml2WMpUPm3
Hf64e3eNUrEwHmyWaK10rG8bVkwtiybbjAcvzg1EQoa1mVsdMG0MrrnCEiES/FmL
dUh/0AoSmiyk21+s022d0TtTD50PQkQYiwdlubF7vj0kVp6wgY2y7sqnQXl1XvRA
pGw5AI26sS2/785vK7k7XbdjENYSa9Fdlg9k6buG0JKQadJzBycBeS8zAFp8Exho
XMaaVNfwIXtDgfMd4agUZtD4WsP/MHoz7YL6XxPQwBBkibWKIHDBF/R0W6IxYR8q
S44JXUDQ7w9yjp6VfBH8ObnyqkEWcioQsdwEZFBb7sj0kevx9qI8Kgxj2btyUF8d
9696DSgl7o6fRPPz/xW2Jo5g8nzFnLx00eVAE5mOMeGbsrGUPub0B7nlL09Lc8bA
Ji/wcOZ8pvhvQB2QhD2nga8LkuVCvjoynwwfy/jvDX8jJ2b2yw4AXaXRpHfgthaU
+0Ld92XlOIOh+5daTxSDNzmpgjQO/ri0ln4tVkcz/o9Ra/Rdn8WvNIHLP+Hp+xtN
BPHDljp31hJKLB5/OyhG5MWwVLayNtzluRLfCpzZD7uPAmvGumcqJVWiHD3+9hao
EhC/ZzZsm3UC7CHqA9ilUE60FgxD1dbF0O+e/I6Ywu2k4cZvXuW7tC9TBHTf9Kg3
gmH1Vz9Cy8NXzRvS9SvvxTbvpu1BR2iHU5QqJcgIBAbkHRSKQcel5EnblMkEV7jr
RTRGaVNjSWJD8H+PehQQH3IILHXrz+YE6TjxTJQAF//QiRRAy3+iHEkxt4jcTplU
KGMykeludWoRSWBJh6wOp2rlzA28cqFsNmUuMSlg7UPGYSAo0FwnmJvgN0zzB+yX
BRN9wvT3bjf47FIdpQtpuXK48Qnrr4/YYEZAkqvMUaHQHjRCkDTLi9RJhttdvFBh
qxdI1uUb4oC2dj0QnxYFgBvcR6oPA6A4Ik+gorqZ01MhKf7xw1wmfymlKs3Rnwmg
NdhQDe4pjin0/m5bmM7hPF51K+1Mq7PREaTQUJ39SRnryoP8E+elhhPnINOdWuUH
IvKmhJiBTEB5/ojCJfekyNDe6Nl54/EGRCkDouaxor9eNfNnAgNTVuHYcAsRZ4hB
lns/T1h1Q3SN73eALbI2oM5PESFRABDoQDlYsQGKmlS9f+s148HJnNzTsDuCEMrP
OZVBh6Pqw9dS7jVY42VCgSW7/ZYiV2FJkepeBBVUfa4Y9sSQDmwhDzNu7j6W8uR1
8aOaiLnJGPw8yjJgM84lIx4ecSDwbeC5lI+Qd8IoMqNJebx+ZuMs1gaYuxK7e3Rc
mMB+qhQii0R4HDdlk/J+A3vz/P2/cSRwqfxANr8uczI73yuXbXroL+wURLqouNgX
OAJfs2i6g2P6kBmLIUWNS/Qc67OUyQIqJrZmM6nOFvN7VU1GGiBLJ4zYfWrWr2Je
jWAGnGuGgOLn6ednYv7JDUmVw7I/W3Y/NX/ZSONRQ6A0DjbYlIj+wfyFUMFCXfX4
xNTNC12pZ6HPh1PMAoyTFX0IWrV4MWBlMAFFF3LDCWBvccXr0jShf330PEndqZLv
3Swjk+jfXxXoojP6/nUnE10RZmAVFgzLyQhQQOgpuCewcncpMdetr8JlLKEW6uYP
4tg0Vt2zm9kMtCJzHs7B6F3tzcJYHqighCJU4RZmbrWsCkFWK9yJ+J5ep3QIWjTX
G8JWAEBM5KSLod5dVCO87pJ4boJra/CpPGLZ3xBFUwGV00FGsnDD5y+7re48TFOP
RHb4o2ZZ7zF2WrY+7fq0PT9+Nvst9R0us88hY6lx9FAs/T05Mu6IWGVtZ/LtSjkz
wqpzfD48rY/V03fBywNXL64MObDQMMDUlS2DQLYZaWPGQebkJknN4F8rcW9Iryun
j6KJdkAMyvwmthHVgARbZzrxMgoBsQcG8M7p3k2rN5362LSUkLmlxagjMxkMd/9C
YIuUPnxV39cElGuRoN+fZNvtAgUE7iAympOZKCfEPgh44096d0SZp2uEOR+FNKYF
JJgku+jF7iWYpxvKJztk5jCWlf7RHHQ+VKKgfRg/pHf5TU4pDDwY8gItzd/s7AFW
2gENIrKB2xVnacIEtBU3jxNcDKzVHhb+7FtgmM+dOxzVg5tU7zF4DUqN2xAK0YiG
lGGVt3hr1pNi4MBlWyaJchscD/NY7aRbA78/XmpKYY7/j6xnS9rZMYeqgs7/8+/E
urshVRxkaxhq+8nsJ2aMrNIMgRZrEuJyeB+d0T+sORAoyl7m8hUCUy/M7G7STpCT
+qeef7VsNonaPg+V/jNuKlcFkPBX0PVXKQ+HbdSGQCZRRRfAXwI+3Z0rs8lfcCw3
Mq9DpSHM/EpRkmfsl8lEfrKtKsskMYlp7o9NDG/XyNYaG2R/sD/0SEHYajl3atwX
YLw9h2jQoZOEcM5n6axw3AHcYb9lQUEl2SnrT7LlOO1Fd6YOQBdj6xTfiIIuvx0q
tz3JU1IcIk6Iv4TJuAhTEoCrqxJXb1Mi08D1UU3yvgKNf1JCtKoA8/rmYEKKiZZn
KJUShnnV8c5swJlULVe0HAHjYBnHboKSu44e0REnuNv68DjNr7rlWU0NpKlH4NXV
Z613sz9ZsLdz8AbNPVdBt0tW2Jq3BRZkTvmFF0kr9laDcgD3rIBaQkmxP2iupW8G
gV8xwBhBiymet+GE4tqoRrzk83omIMrgfmUbHh51eHDCqMnGx4jLU+MWjmCC9qii
csN0ag0bEVALRe30o9ntU9LmLoBZBmam+q/bFIf+LvG7M2jTczlxdjI0MdA8mlBy
7K14Znax6O3yJvjicusofeJedy4OkXyXO+BYBlqfBFW9xPsDSQjwbNGrLw7M3MP9
Ei0YmlSLW9LBze8ubYkMvjYnMQjzfPh7kNFLS9TlT1VQWvdZxm+/hKRoXPjXH1fi
oDGt+QySD/lrnQdS1qPiijVIsvXgB65qw3P4ymONJI4N/87g4hBGnBNAOrrLa9BE
6kA0fbZOVFSuL0+4XV6XOXAW8jsNw0i85Y273ryVNybPinHKfdsdx30Zr6L68tY0
Gk1m5pJ/Hh5LWJtoaYAKirIiqlVfeWc0e9Vzwn07flx61NauGLfJ6zts2jtQhSXF
NamXVhP/t2Wj91UNFGAB6BlKkZwRf7XcdbFqZy8Fb3JxQguxSaFaU3ayFQFJdCuP
89m3zIUmIjNjzRZ/TUY1JsN6NtHjzswqTNgsqj/01f0JXayHeVej4GW5xqJFCziY
OL7SUfu2SigDEuISE+wxhLqNRC1P0LQHT01McWk9Aq/T7C+hLonI6EP/IWxTEzJM
NZdAdspC+I00oI0j2ONklmPR3K/YeHWqM/iegeF38eF7TGpxC2nBQXUgtXFKuyiy
/K6UXqeanLSVHZSIHLj+hCe/BB0PyXYvwmV1D2zTfusMbOYY5u1WO41gKjmeYLRO
dkD9V+vMDTvwyU+ESywTSnO4EyUzu2Wx0Dv3iqn44uySS0F8oAWmmV9ZQu0pQhxY
7egmF5qy7yCM8Xp79MZ49quSYMeX6mRkblGzlYWq1iGEY1l7zoHMSGYk4xbeRzTP
wCBqbY2iNBDy9l35UdxVe7chbfM1CKyMli5By8RVLebC1ljPJJwvENf7q1vsbsZ8
XapeSw9NqDTSAvSude6K5A1Z599ae8+BnTdHzROtliSDL4qHolPoBD3UgFysND38
Y3MCjq6N03oT4mcuUFFLsbk0wDh8+mVuyQfADq5Q3OQSfmIN8UqJbXfxjfBTA+o8
/NzI44vxTd/h3AAitiCnaNG+KQIUrhIINTvj42/1Aly7xxvtldnBgC9jHZxiFsH0
kNU9W2ByM6iZDwwq6rmWT0Q3HQeLbQvm1PeIJ0IEz8CQDfz16wi6tzxZ7nAPG1mM
yoOMmdHv5Qgkbcqj3+8oUpAlB00+KIqS8X/y16FGE5gou/AGqT4GLrVKORHi/fdp
vxdP8dnVa241b5EDAZwgTIzoT16Y0z/AaEe0s+zJB7IQFVVoLCglbUK0bgGNp8/c
PpzRhvD/52U7L5i+H7bAlmKU+18S8o2760eQq2K3uUdwl9zuuHGptgbFfxPQSFXE
qPNNbAdtRbOstxyG+Ti57NpgNqTxeFs+DBX4eKY6N+f6TQGYn6UbCJkWsjjIwq3Q
83qSMNe0z9dzu/DWjqnfdPr1GuCvzr+YhTmO3/A26D+7EkzKXSj4N81uCstD5tXP
mdYUSNwTlKDcNgzHj9oSNHbkJeB1+JdAmRMTrf4ADuqxv5T7OerZIxI2yZeFOTh8
k2OHq6nEprmENpT7OU1vjbkXIKV44iJDErZBNWp5r9BxH4oA9IX+EbWLlf1FsIs+
x/xqT0KbddmDuzwqv3ZNdWRlcRY0/S36ZzfWEECvV/m+KOT9R/4fTChIKJg4+pyA
PiPKqdLp+veQ7s9+tMQKQXDMHyRj2EBZvkKG8iMcfL7M5kdfge2v8idVN4iY6bPB
UprwH4Sk2M9unJHP+LmSyjM/4Un7wS3akyrv94+OXxf0WZ+tcu3CaaPNdPAgJlQc
XuCDXTUPR1dfIMeV4JIMDz6s554PES9rgpmtqT0cE7w9IZ5/n2irH01wTUFPv7Ey
v+SUMp+mxoOHPbfO7xbTEbN702lwXrEnyT/wML+aCzc2LYfPfKpvzF6rmfMzkWNu
f8OSNT2ggFF/eFiRKld8S5oAPVGtGpxN2gkeCrL8YqecswWO0feaVNNmzNdisgSE
ikLTGtxlZDIXVGuhfSfha22V+L7BhIOLRX0joUQuaiYnCHpzy9TPvF4ySKJAUUEM
xenfzKC175OtxYJdfOkC2yW8Wb2Y9gjhYDRorWyHsa6a7VYjKfhfPDbmxbJc4oSH
XJp/oyOvA41jLdcQy6wBYJhOnFt4Cm/VT0XVn/WYOR7G7vtZiCcXIXE4AK8WzJz6
tLUZzjc+MP3Mm/KhW5berdnZeQ42degid91+zwqSvNzdndc0Z/sNJjEHacfazz5d
0veU25D2QkQV1rqrP6k5OXgbDbxHOO/9C1ZV01xjyW8VGCJFAYp2CISIVjEjgJ4p
H8NlD60AfUtU4gcq+V72YBdhTZHv4XmlWsK/xfI1I5bcz0pDKLACu/f98fyY98vc
axboK3JvV58iToY9FWLtUweZlTg7HxcXMSdzB/R+lBXOaYrPJytDvaGDNpjX/Oz1
M0px/MY5r3GFFetPTPkNfo2dnFWeOxiZ7plc9jhN0JqNkyDqETq8+sy6h/+63vNJ
uRe5TrocTdDdZPx+yUfYW0606/x1CNL960w0+G/KuzgAbijzYnFRSi64gNNlAtgc
Js+WT05gF6mu8fv8zt1kX5XQ/xQO40oNM3oaPJIOaEd7Pkm3UdwddcLOL0INWOL8
QBFAwk+KVEoXr/3N3jhd/Q3GAQrkDeKHlOX1/vMo3ro/hPt1e3yn5dWcX0f/v8fg
mLRPT7wyC+nkmrJvardsUovxPH9moiCxWBdu/J+XDRz6SVetVtBh3aVo34JGnHew
YbdXfSpJ2TW4zEbzIufSj7eSO8EmKqoaO6Ni2flA9GpqAvony13WDK4tZsb0fPqJ
+xvlWyXJAgcUDbBvyPkduJKugu9a961G5JpdmfJBBOvYsd72IgjhBQPxY/Pv6x/W
seRvN5FzALXeCQtFFRuhhWDLaMNMU2CNrKHt9QyD9OkkHDIJ5O6Wjc4A+WgfJNbL
SpPU+38LDJNMjX7h7fuEq0PXh2lcPpq5IjAvt7nV76QIH1duYgl7146nFh8XYWiQ
9UPW9Is+qwx7qVtDYTXaPXXNpAEX+a9OAGL76RuqLs8hW0OrqyrlZ7HUDflwaIPl
wwmiCZ4ZmllI8XC/KWGdi7putEOG1sDVZiT4uGxrdN4pOWFiAKNo8NQ1qbQQyojo
QNIc9oL2PiswgOax6as7sjL6JAeRFB1q8pJb+MqVDEU4G2DufQQ4DHbGJmXkgpos
gcMB6gUcMl8y3GFz8D/+AvJq4aau6LQbZHtZ6G2TTb+pDXvFwDlhG6/SQUgHgSBL
AMk3U/fASnHbbDQT5TmuzmHsZRCGEIo567x295SOaSCG1Od7xcYPp2clLBfIjX1c
5tVsYjSYw0YieqNwWULHWt1HeLHIE3ftzr3JE+fEimaWbDqoo6QKQxWv9fpjZhvr
d6STnqA9wlWQUuxDDwX9xFQFL8/FhU05SHgjmApBa1UwnKKpREXHswxP7p8mIGAb
dVjGJZUXwjUjFiBxb4DZovZV7o/rXUALH3C30paRe728rag01kNqjNYtcI0twTRW
JVkPCtIVjXZJPTvb6RdHpMODY73GY4kTxcDGgtcFCDAgrU2kUUBoIaI266NOY8kW
eMRg5GxPYnd2F6Btq/UqpwnYAor12Ev/3uYn+6Kjl0ggD1ET5lKqnsFtC9RWRZF4
b3aeaFIUpGvFnTrwGxMtnA5irrtegnHbQmgw6c3jaKzy21HOk30qQbqhpPca6aJO
JtyzCHViLW6Jh5J3+i9gMB4oV04rpvVAp3PQrrLHXEn6sYfAYGVOT94g5lltLqdY
0+g4qGOO95Y5YHM7oXbIHFNS+xVnps9Mr1fdj3Yby9i2JfNlem4hevPqjzRVNv+Z
Jv0MLJQwoi6QqjURubQD20uMJ2KUxQCxAgQgVTdz+cYuUPel11yOSxV4dfa0NnCh
qOTyqaFayBg+XgvB2OnuBGbHtHfBENdRoEn5V4R/t20kgDuwqMCNnL/CnnbIFC02
+cfYke+3UbSrcsz+MEUY5xAWCcWPx8iLBTvlooa6yN+6WkxeIBRxa+Y7pdIbNB5j
mXEnnUeuWq2T+He8cyY/q2qS6TmhuYPdC+9wiWir+cP2LpRJl0n7aYfOg+3d+12L
mgEphABeXW97LQemKRXPjKvhXsbxdwzydLU0YoQbJLcg8T1MmEisTByOJiMvZ1pQ
MYPNGMXCsip8VpbgdtV+E6HyfgwMu9T9W72qnRLhUtG886mX6onSPmYgwqQQ2Nke
2DEk8KWk844AT/tIzJoDM3zBjZ10z/1IKDVLCgMA/0sF9OU788aYhdCFptyxx6Kg
oEQxQeZPha0H+DEduy7G8H0RLx4kqjQluTtnhkoezI8gavPwmYsUhhJ/Q/0pK2vQ
7hOrzExYZxWBx08ph7eaX/Pb3UOVgs2gl2RjwMTH3o4AKPOoGBOSGRhMMK627uPW
IkqkIbsVGqOEAQPkrb4qTunZisXepE91bK9m+c5Z/RHHpePLYea3oy6Fx3Z22xKg
IyNOin/7Vv+o78zB84VDb685Ir1W3HorUdNWRKZLYuIeYstPEVJ62leP2j48uL6d
tNkGCOcE+TFJcxBLQZFPoJMybBt6FgbQQiCksqg2dPgrAgkYX8WlgcnIOIX3QjsO
0/8QY/NjLtLZJjyfKHFEvzbyJydpxAVajJL8F89dbe0aSyjwTUIXPJdKdRSlOQD/
Vm+8xcMzezQMkArVlmkgUb6l7Om+z5CQqCa8mZm/1Ke1t85pNsbU1wHoHEBhsoTQ
ZaQIKbP81o58v+/gu/lRUAa6GQmC909MOt5aVblcViaT8sbbgzBpOdTyW4v+DFQA
Fk/DT5XtpYPHK6fZStAg0kxCuSUiXisw7plsg0kpG+lkJ99tbDEh12s/5itbXFXl
uPFGq/17Td6hY/kt9pQF+motFNmaj3dq9d6ya2IsnBFjrOXLoxtsytxzwfJTtJ7e
V++71Eamy+zkLkVLpH8TpJJCQ4OQ4Kx0Fq/x9/GjJzi4UWdcbcUx7q2vEFvqgG/p
l+JbR/p64OtIXLqjqc7xPBcxFe9vwTjKzsHH0PJuRPTX1OAwOhjs8cHaeTixvnzW
DiORTjtgvVNoE5AFy/fBlbHBbZqoNWeiJMjl8XNRAr3TSzX2nmBK3imKrC4sWYdS
gRWgdhe2IN1RR2JtagYWYHlWrJe2eMSyweP6MvFxYHPS/EGATO9aYkg+ViMrwBEx
FssC0p2znL0/pHnW+JONdSFaPYIuft/tq8SgVbCK9pvmFWDvKxqYp5xOlAp9idvq
P454dlpqCQbPSO3XzUfq/D3d0W5teAs+ts8DPdhXhd18687BOLHfZCJpFrMxe0tk
ObNog/Hv6n9QkZlyCuYW1xW7jpRi/3ZTXEMExOMusyYrvdVTN3Ip3Cb8NVDhsSp3
4sRVljy5hb2MFZSAaVvDIAJubIEhn7rgJQbqGGmLo4knr8jdBZckkD0wP4h+txyn
aUHqjWh6VrCCoduGR8zDdHHkkQ3qGEXPB1RLJrqOem99be61v77vAPgx3QSKzsbf
vfI1b5l0/dNvfP21Zn9Vyah/YYDxzPFLrd9OLtYXWg2BZ1t+AY2mVxv0Dk6RYrPc
CIMSOFRfOrWvMEWeowdyJpJoLpz+6O8R7dgGCkoE287wyka5rpmgz0Yv+XnEdxgR
jaaeI+idCDszVSL6RyAvOyNIMNa5BpmOJswqSiGw8gze1xyHbikHDBLVOLPdun1o
DoIMPav+vp2xg71Grb+Oduksa3rvUnm6FByd6SEIg+mVfmj6kvhzoPfLThCOeFss
WGaJ5k5z0tFta5WIc4UwgZYyqZ+F0ERRgfLxgE5woglabjAdRvGPiEGk8B43w59w
/Rr01aSVmVviJhYv4zwtfwagFJN71SgZaNgZMGNzimJZ413AyEjBfufu3fASwshL
LjAREhWsxBIJJxr4xjyYNDhOFirudkA+ohWQ+Ic6S8wAO5IC9XiOeFlGKt/ScCf3
jEorZ0bR8Akm73z7pT+ytzUXBl93szbQ9Mn5eHCsZggh7ZHNLnI/V+luhpfr7IKJ
/N623JB9fHSHs7s8pUvQI6FQXvO0xuEw1HUZHZqvW2a7C7j5E78oPLEvfV0U/sm9
GtmiQUES7JNCPbQcBAglnEUZgx4HLXzsxd6ZdAVtJ+U7Lrf3zFG5ASDcQsJNhfeT
7E1KB7kK0ubSVekrJs7XZkiwQMWRWsN3SUoBpAT+/BvaE1VVmIXAfEcbpsOtHi14
N2pl22gYFFArr4QRfyKQpAIZd08AvteFtnidhK9xM6E/9Ybxo4zX4fvB8qyyis9h
4/9fkpJDXuFmKFDJ1+mMmhvLg5eNjn3kC/7wd7DKALSI5kY5brLDBbQt+gwF1wqn
uDy5SLAQeDUfBSzvBE3iAfLkWIIfmZIhuUnVHPLG3b9UNLyOG7YldkG0Hk6YKJHb
hIE5YohFYoSX2PWRNMgXb+EmGSirlkjnFuntsz05O84Gf31jefu6LjvOglfgEKl7
HLKYMx3Z3U3xH5jFwMg2ttnzi7lgAppFJjOYl8oxZD7H4QJCY2CpLFh2EejznuEH
uxQJH1ttQd14RP5mwNHlQ+24aGYX0bCHBU/iTjLRjBA1rqEDva/YWHPLkPY0O5dS
Nke3F+Pde7kIgHolgFpTIiVrqOozy97/oJg3poPNUIyLJysLnUNxZu5Y2MzkuHFW
HW5KOiZrvFglzXJyWBjvNdRxBLilbd2QaYSZVwsHQ0AROQwj3Fz+sCCT2jl4JGUl
T3QmhbHru2Qd2cqIJ0s5A97Y4+8RCJib3AVRGExWAg0bjR1bk5k7+EWgYUKsq/5B
7ZyvO8OtmYbB0JIuZ+52lRRJEE2Yi9Z0maJ9MMw31JWH4B9JlUIfeeu6kzxIPIXv
JkMzpLWNIissrqvqTB3lJmADt+JLkOkIJeq1m4BTkuRvfRqSJ/gEwMgglZPUyHvW
MIQkyC86rdBI+zR4Sgmw3JSYNHdFL7YA4uzvhcy3DrkR0GpZgkLin8PkVbg+AnN9
fznQRqbDl0sIU1Zx7d6k/11Wt5ZU8UoB3Tx773stFLnRfADHC8/MmDMFYxdAS4VZ
NFaBicdYtDPsBRb4wPFjpAdnXbMVf1KSTGrp37O84ZOAbKDFindDuEfxSGTIJubL
Pxz8jzJSykNjD01mbL+mHUOdaLl1qXbVU/LrcTrei7snhKs+XaXosz5FS6qhbkgf
dK4G95WbGZ/3s3KO4axf7Lm2/cM97xMxD6yH+jln7QKl9VhN1RC4TvhblGBtzbq8
jg2t6Sw/CsbW9v0MXlJTKWrjNti0cDE0Y5cJNW8aADrVR7v/cbVSbojJ508TNP0c
sAFBsOcMNUZZ0MErzqf6GodC2Adz6Gt5/xfXDcPBQE9XJQL/QCEMnstBRQGAJGjy
s/t3E0TzcZZkYvRJUoF6tXL3nYPRvkjwpAfb9ZeUJJ0XoxoODFiiU/NxpKLCgOqM
L8ZtXv4AjMmAgZnCXNt4iMGhLv+HadlGgw1FH0I/AO1P3mBE/Vv1kOnWdKhVDInU
eoz5FS5Oj5RalqXEkEP+XJKUYghCMc4t/zeQTRd3vpHv++oUkM+VzODY3Ja9pZCu
rv5TAf51388JDbjEFS2uwrVCOZhKu7z91Z9b0N3MfaqiuuUgp95RkugFgvHTDK1C
dCT2G/nPmgxKgSKVWPvEcKxaz5157v+3HzxEP8kXUOucrYSUhSREMVWiRPDK/QHZ
Y+QleXRMKVI2RjeYDEEA5FbPMSQsbDf7liR1+TRZ4lOoUZTexp1W3HGaqDziDwFK
+zPagA2nI+XaHVlnWDq0SM7Hl619rUB6AcqPr6Df43fx+i2lrN5WVppmbKpaLm3R
3KHw/9JYhtaSf1kuy2YxQQeEtKHd2GvzXDXmwTlUpe8RUuI4vlAgA9TaFt2hZCGc
DYw3Vz1rG54nS0Cnj2UGuPsSRqVH8LImSuMLg9bqcrixrV/b0nyxlGt90yhPFgaL
4wDMKt4oKT7UqTWEZ8fDdgAIdculPB+lA5KtNY0ZgAIC8Jondbhio2vd9d8fRzLq
bTNm790yQIKzpPYI4br2gvdKOwDiquMBQRS6GhV9QEcCAB/1T8yPSp6paR6rgSPL
flBoFk3C8XW7jtmLVSJ4rVHYQH4bxyXJVSpP3FbVI2t+RwzXdpwhf5fbwACkmZPE
j3glHG+xbpv8Qm+IgOyFCREyYJpRMlMiQyJfCjWzsgtpKhxtbsZXEOx17816b831
gV/tv8atC5vf3Mc/dQHFVN+9+LDuDUa3QdN1VOovKR2xPlYu8TjwZSbuhUBt5eAc
+Iy2p/JkNFR/Vj6fnZ+no4n+Iof4vst0bXdR6Xf9gTRV47VzyclF6aHR17HYpyr4
mhjrnTmPL2azavHvQeRf6ajxTsefjdHYO+nO0TmixfVjpIMxNzS772N15/1/tChC
vXPa/5fPDU8XRoDIJ0RbbWG0l1tmLZIVIZ6AqHO+Z0knohHchMt7HecMP0xGjLYd
Ua+DyIPAUeRSAZ7FwSb7ryePjVDR1RKmYZpLMdEkvGAM9vp2FXjFATRIOtQ8byRm
qzqMSqqUXySilOu60U3mdFdQpBdJx8/t9sY3n8mEI7G0Rq8ithihJSsfrqkTJ6fL
pcRIwqQ23o/tdnUKRqJyPw7aLpEeSEVmvQ5XlkFtemcw6zvQ5qgkiQ4usmE0cRLt
0CTlBn8N/gbIIw0guB+o6EMpibc6vbglbgdeS3r+uVAhpAqxfTAc68NmwsjjVDh7
ZeP+2Gn/RKfgt14MR1yfM+qaTdsEaXGgP+LUD6d0GfM7+hzEz5V+eJITvOeUVy7p
r8jtSsS5WpyYLJ0oafm2cODcE2i5WeW+CHrgf5q+ZI0VhAUNgXWfjd77nQosYyGd
oFlc69dxWRrpyx+hgYYjo1vIEsrvBJxMgqkZylQSB0nxfpdrbwdpysXOrKAgysNE
QicQHX/2tL0SDVQX7lb0ajF9WiyWzuSNpxhO4rxN4EeW2wsYJCk0E44jNVafei7K
2acYcwrqyAHcRN/w/OFCDTkL55pMR8hJY5Iu/Jt3D2LoTBncO7395TYsMXzb9ENf
pgPSlvpTyiyeYkWrgDgkI8gpPDQZ9u2w5Syhgp4MV+6JcF/f+vhOxtzC/urTRbSt
Oj5xub+FJbZMHvZKnMdRq3gfd9HsFzgtXdU7v9mWE2Czyg/4T2kangeNGY2azmGs
syRtcS2ydibCy9ubGgsOLD6cyqpkY5hlvevKSw9A5wMLEbvuRl1v56WPO+wrRb6l
rYfTuTvTDYuoUkUtu7UuMXYfBcR+Soj3rDZkABFebJi/teQbi6yrTrMjXObFpfIw
P0DW9BIEtJS6nx4xV0ivm6Qsbv+aUYqkDKAuedYXXRMAjuZIPJLHYqfbcdG7uRm6
/TKQuYnFM9mXA+DH3/nVMOKlINwyLffnXRkkvZaYLEnCtimgjKrj2N/aQ5dT8KyN
okKZ3jg/jlUdltV8KW8GpMQ+pxzLAkguYDHRWZUuLHCTIWgxfhMmHD2ZzkpjOGne
59E+MZr5ll9qu9aD8GLGAyWsvBB+vyI0yVeHz61ObDsB+y+lbIfjqjIOfLY6B8H2
8Ivuo1S37kDNdpn+XKApt3XKcmm3OaTptR6wu82fNDADoN83LxTB5iANQWVhfRnH
9T65ObCRvb5iDnXrXykdt8zHpIfSzGjr7W5AA3lLmNKrE5eNvv/czsQ7A+Modibo
z4eKWqUda37C6jgCx/WZtUk02MIsNmw2GNKH6tHS/hgYDAsvREMzvVXQpmYYPKVe
pzg8GlHDhpnF4cO1ns+6v9RRXsA6TLcPdy5I6s8B9HVXaNKMCST9jYT3jfzlvw62
nA6JLETOTfYLTlb+U2CoqypriH5nd6TgFsefDuJMKVdK/tccC1uScs1MJhqjfjF8
Qb8kCkRFRSB0+88Z8iNRWEDj/nQLnUt0k/aBpQlp7McKmrDbMDg7GaiboCkrEW1L
4Y1wieBcgWOi/hmB8xWNqhZadObK4Sv6/cvX4aJh3C12EuQZyyz/KIIxH6HBf9Tv
0fsJBw1llLRedtTAkrm9/oIhzEYD+dzfuFDFMqbORqGF6Js1N6KnQHjxxWNOG2Su
z+W1DBu3GGe1LcecXqVP/su2Hp5jddFS1QnkgA2CK+CHa1CmHxh01XQ18rknHPkP
PKNmO8WOfvG2yckBDl4vvde4nhQRy4l/Ikfp0g9MZTTm3nHxlxSPpQSK587JVCe0
rVyIRDL0J8zxslUsgXZMX3EHp+TQqDFf01Ha8je4ezk996u2hwoVjMD5pViRpNgF
V9xd1DX5yijbOJfWq4UhW59EeY9ycLyOuyDmgsPIPDCCvJRCkymVunJ1/5Vi5Y0Y
scHRPDewf3kLfAMhKamYtOJ6RMHch4zBCyLixpjXEKTJ7m6AO7Fq5m6um2WWzDD/
h9MZJm+6/wOIeVd5YnDYh6G/2+QE0/9ycgacGbjuEKytq/8JIcVl0De/EJH+RiX5
nC6ya6V0dc6zQLbd7hPAo1noBMELi03Hc2roqGuWQGfRYvg8kZnV8PwsqW+Pq4zC
t3k6RrP4JcCIpkcR/m+NIvEyUp4WCab+Ypn7xVjDpgFxvw7xagi2paGQPT2q05n6
JSg7h2ghADUp/x0edmkD/EZpQDQCgsPymV6UYGNBL9LmNMv+5OJuUTVfaMLwOOhq
7e9UUBXmbzvHqqOjulhJroRzf7xfhd7JPvtwPjwNfReg3mkz6mxS1WfqS4GvP+Z7
8co7LmDOjJGEmYGi5S4OsUju45GBgXSWKH3p1r5A0RkEYAF6jGo++iT0wEguchVe
WNle4Zp8K52FSdOIFozWVLoYoHria6Vx5ta7r2ivOnwDF6870WB8yerMRnAfbYH8
JtFqUi0IkAivrWH+zarZ3HoO2xuoBuf3M9qBGfB03n6VicqyZ+h1KzjNU2KUtM2e
FKMYQS42CrBZ9Hgz20tzsrU9idRmTXpYpM1A9dW19RgnGLUAKLFsgt+jCB7nNHwf
BQpYAIKF6Y4/olBsbNVEZspifdeSFTGUtSG94+d5CfipeRW0vfBw/vCnpHWgX2ch
zHbdDH/VbbFJYPTLrpAd/fOW8JLv992qkiK1a2pbGuUf1zMofb1kqCClNwASfv52
5oiSGgtHo/Gk7DekQSd9qBXKzNypl6lDWeJbl3IiIF7GqzP02nucy0Js9tNUVC6W
Tcp4fXpRdNbw/9PZxcRIem5GzhcXzbkRdneUB08oilTCi/ZXCy1pC3t5Wq3/nM6j
dSGaWAD45aECGRDsDg36lkST2y++W6/1SQaJ+baVn/tJy0+T/URzZpAXKvCJtk1j
H1yOSIqPLiUY7qvvPa3tcrMqQQw6/h18DRy7yVr58B+rVZt9ZMF6/pkCmB92CMyg
QLYuy/neA2JgZHWN0x7bZ3JA3sU1ru85y3T5nXqbs62spfmOAcauGk21u8pJH7Nc
9J1LFFyFfVBErKHVgXu9lXhCgQKfeEaXcERkrPoaSYrNuxBVO9n9WWQ07KKdmZlv
Ibegy086vFWGfKW56sVc17WWXzB8ebfSvKm9J2oxT+w0NaRF0XLQ0VhQCPe4p7sb
Ih3y+4brWaeJUxPyZXs1D/ZBXIfXEPRw4B6VsBZdvYBjYxHMkH7V45AX/T1gSP5g
+osVOAC+c93WI1YALGZ5Ms1lFGWGmribBDLwE51wry5jcLfAAnzgUZsg+gL1kL3a
yKl4okhNjrKNRFCOqpdcJke5DHY8fGi3fanGmbz3fqy3D7NnqU3iaV79wyFvgJp5
P6uDWDIV7Ls0Y3VZw1GG0Mf28gpYAjLrbQeAz7slt23gzd70/TNCE7ou4eKfqD7C
nkmxs/yCKGVVNGJ9PK/xVxgZdiPSZbGd0wCTX59vGOHXnbUZ3VF0dZwRu7sk6Z73
80RSu/SEvw1s03lMPguiq3Jc5Z1tMkAlYPGjqmLuRQuymPv8w6Z6wxd1v85E9ahJ
V10Xm5tUz4VvwvHMc+w9hAldmmIX3hSPsJLiqICtC8Zkk33kbolWs1t3Sksm+51X
N+Zd9TUdSlvEuv9rMyhXNuOx+HZjEdI8mfEL4SNHrFdx+UPw3orOMReg/IdHzGyv
9n5ILfHeTodbEEwhDWC69+Tu8ZjOeoc80pnNfhs3jXbN8feIP7T/daaN1/lX6+Yx
glNv6t4FoT2w6J1+iq8JXdQqEbjycw3e5dY22ZGDWdGDo8dVc6sQajd2Bio1AiQA
IUSEPk3zuatAwKDTjOyu8vvs0gwUoYLwDUbu4Af7twYOvLjNiZch/rbRPlkTBMSW
bisUmxnymAY3jculMWTjuLjdfhnnBEu4O9kLXcEcp2lYb6+4O/hgi8vcnVmPU/Oz
qBX2zKqk0YmFCx3bIVkEOKlJP/UQVyXIp7T24AvT6vPzNDiI8zpXTfHsMaO2SIar
m5gBoJGHKGHoBwuO8zBwmmfqDi1JLhB+K/XKwUaoAcsb+aZZQpR6hiYUxDki9FWk
SLVmrCuzVJ18pQ/XxPNMZ/Br2Bk6PMyCFWJDRNRrtgLCxcLeEzxmNlG11VxqVNiX
ZfmeGkh7j5Hqjq6k1VvlG0jismtB1IktlfCQZzEcuGJduOxLbSfXBwQ5mwyYm00I
dz+4Qd5GgHR1ZrLxTwy4cikYFMy/iMyNldqN32y1JACiLUszmq1IJ4IqSWQlUOD2
ILAj+ew0wGSaoogNr7hWDkKW1ATcCVixhfKEau65TLYjtBAGV23hafBIzXHhATiB
RdkoDfO9UycPaBJy0bg84R3ouNGTJRVS9Zj9VTRa7JZxHxJhMMq4zUFS0+ZjWmvZ
cMyawOYtbTTEGn38UH/yxNZ4LRqol/80zZSTPBuL4KW0gn6K5ABSbcVLWo2giDtw
J63Tu+HoEq1v2k6ym/3ixJBNydAHICN5TUaA12zReq6TmSRlWDIxhretxYJNPqkc
HGpEqiu6Iqt5QDK12VS64DTgYik58lzkauKNzVuFX7xqiO2njTH9wKaoIagSgpYf
eb/LtgeYoN0BFHiiD2rRwasZY71YPwoLm1GjzuCPYIc63qvTI920d/YMpAQGjp1D
DPXZJz4A+FfPsCjZfPoAh5UTQbMmFfPEkY/WtiD4LswLd4kxem7Nni9JnZwGX0CN
KSKoNqSlg8YghviYt73k6haQhI6kHuOGjErQ6EZGow0GYVBhWtatoGE5TqZmxfnQ
ET2vxtexjpFi5EmQvBeD8+7OSa5/3D58PYNKimQ7Rf2b7OysYbiGc5PQID5GvIkw
PPb2WCXeUq7NdK1ELcsmF80z51/FDMhdUVDLU84CePWf/FZbUhveGR9wcBE+Hc22
HthTkv86m1XrVaghLKKdWSL1g+rJ2lfwSvD/ajg4dRrSgccd3ObkXH7BNWhErEKg
2MYYGzRiXv5pf7OqOH+pWSgKzLMszk77HAu1sQ5bzwWSCijP2qgpg98UIpTDbd2k
W6+61cY5482a/zpORJtE9gBrAQsD/TM5wkHXG4JSqXedc7JDycent2a3hWGiJcZV
zKY+oXmeq3XHwnoTcU2Mx2+vdQspwUcoXVds/eeKYMhLXU6FYNUigaIKr49qU85S
45C865PIz1tUg4niFyNb0SoMDFeg/5pDYo9Bua2bE7ITiZQ4jNs6SkVv7s94Fzeo
4pHBTO4asffOA8H52osbgkimb+sibZTdzxt6N5Wwj83Il5iDx5nEgq0p9y44gakC
fi3ZFfelG5KwQQ9Jt2EozoSQqQxTUJF7awDGAabxVXurnJ5WjmTazMqiJJ2fucQX
CqvZ+5ohtqUhzBYaDCaRLC/TZYkA+63yfDZ1quMHZd7kIJ7T+XYqk31GvN2wb3Sb
fO7VbHqlZ763bF0B0bp0m+yLnSYjO4soy9auIZ6PBjqcqGCFEsgSjujN4RhsacNT
u7WCvtdEE4XVaVyIW3q7uZ2WkXGtSwKh3vAk0tYSuXd8STsC2fffuEF5saiSVgQI
tsFcHiX/MAyOKA2VMreVNfv+usOoDAg2g2ehF1pInRVjIqWuKKlcBMxeSKHI61pf
xlbTeSWm4nNc2pFaQsSEMdkxMIh9dIzdRPBh7TvlTvEkaDO0Z3HJp3ISs9sxSOp2
+M6rzL93nZoTaV6vGXTKvE8h3nyvRqhcb+gob3keheEamSTcAAyEBPKlCwycI0e2
Xu1TV7NVJ3mmBDL3/K7pEKasN+YeNA9KmFeH620s33aeCG/qCL2Sd+Dx0mY/w3iE
W8bl9XcuLHgw7fYbmRmiqw9v8tY0+ld7LFIc6reFzFj1a2r655Gip6ZSg8QrPhAj
XyMaBFN9EL8ans7ni6JHKHLo0cIjUTXNoNT1hn9VjCpyDp533RwrjkxtRhBfjCU3
zn086emIwb6CU3phNRZdH+2MiIvrxQHVrJcfUyXCpckQD/58K4nLOveyjQeJWxOQ
yVbe7DRGFWFP5PJchHhyhRQ0jyyco2zzGafGLyMD8k5O+YtEzM7oJvOicYaLbmae
wVLbSbdExin03ItsSoXJd1AkV11OyXu/rJnGLREi2FuTH3sk12ECvIww1kAoqTwC
crozRmAWIqIfm8056kSWRMSZXCksmaLxQJ1wzSJDsiXZuXbeU5VIv833riXGdIW+
ow2oXeADZHJ4vqAX/HPK/Kc/HKY4YLOGrdj57MFXaomxH02y0tilsVPv94UmvqqB
b49Ub4DmGNBmrxSNwYOVWE6uTiEQD7qpIZuG/zxYG0RgMVG6BEvnMFzxJZ8r9Vmd
uc7ZB12x5EtFO/J+gcP8gMa7JizpkESEitP7W7KdpxFqRwf+8BMPWsYlhvJj9Md/
vqY09tO1dB9MWDvEK/mW72QevCx9HV8n/d5XZiFrewybMxTPOS23GnLPzbwJXIkF
PoIN+LH0fl0aWLdY/3oczuxFay7bZL8Igxc4p234yGnRg2qrzpPMlHwkPAjTSRcZ
M1DHvT4lbPYYkjyBfSNCqZziUJxMGLJNDfqrlnJgYeP+eo+nhRRmdc1Jcp+rqoqb
+5qZVpcUxPbpegag/0bCVM2JQnfJDzy7rfKw62XdwS4hZr8S/C9TJMXplbI7SKhI
iq2E1vPAUjxgyf1Ve3PsRT9hwDIGhhewMqIMc+CGir4YqcWXY4diJrUKsvVsvyLX
ttEmLR+ChWP43mWGv498j9SBEfgSgEAPsVCC3hB2R+q7iQq1RsmojIgOhm/d1qP1
OZStT+dvQ8vwA0Q+MXDaHcdDiXPQi3OfexjDYGzM0+BkrScBUmstMBQtoo8akqUo
tYu+mMzKh+KlO4RtVS4ryWTmnqEbgdSkWZ6QRtDxoh6T2P2Jjm9LuLtqvGfNf7vR
4a20288eRPkOk0N0rPnrumHBaTXjlnOEihzv+BkdTNcZoO3zvG46JF6O5d2ZSusB
+eRQKy37O3M8QkP0HYOOySSlCQFn/l/FpJrcgG0DSB7AkhXlyuCyge8uWiQjQFUd
V4o5BybejBqL/UcA140u6uFIJ/EMQmV5C11sHyEl35VfSSHa2y9bvePBs+UBpMU1
fBGz5ZqKQ+vBcifdUR53aSM6BFVmdG2X0zmax/wOnhxhWXM7bJbxLRXyR8mE28CD
SZUTGKTCib6v79ZXSBN+72quYthkWkrKViWcutjaIs3bBDQZPGoeZ1F4GbGwBbwf
IcH3Kx4VhjbrDjVOgjuat4f6Dpg5HOdZYwsa6JRp2nOud6hh7Z8me7+Q6VPMejCM
C32LGY2azZap6lBnJtNgPk8vQNidJQENCq/PnDraqDN4ghLvtwDNKlZKzlJU7Qad
vm9WYzpVXhNkuBwYHUEuKmyS2Rka97XXXoTDwQukKfVJzihb0jQd+OGBCls3xKDa
2i2Va5S9rg+z3ClikEDvgcs1bfomAsvnPrBLwVKdTcEvTXBCNyTsWflBgaMddSE0
4UafiS7Pe2NFKcQCZxqgLKyfSJ1F4INKu7eF/rH4FWED/Yhal56Q3a8ZshbMBJNP
TyPC2S1Mo4wLU5qi7xlCHeMUgVC52XaJ7xJYcTTGxpTylsOrw6z8VfbkXzxWLnuB
Pj7TvieOLQpPoCcTADFpMn28OC/1Pf3oNyDrhqNYd0P6B/PAbKPfizaYyrCHwYPb
76b1qv+goeMG8QZQ0PYQCSovd+IQ3fZF2nuXSJv/f0I6DyQbUztaq9OsKf1cURop
YUBT5VLMoBySl8nTos74yBO6xW7siuVfi6lJn1RLOtB/Y04+t1mWNr8ymc3vN04J
roIH8VHHSLhOAdtG85cjq+vPTQt/BbbiKIGz5Tlmfg95Xb96HEfsi1thX8WJHUNt
gznL5DUpLKaIApI9KKYxMvVrvNuD3RZ0EtOLLA0BDoGJIGshVVWmFlGq73bwF1xa
spG6r+qU4G0COlxJDZAeIzMw9uaU9Z7OREqw37juP00Xk6kDNQ8V/uySsbAHip72
QhYkHsI4ylpF/3cw4yI1Bfq5dqn62AwqeicUPP1zUf09YPqaNO6N9HzWiPdTuXdV
MI9MV9MeUYFBntmXlg9HFms/T/uOg+nm+5WDcIZ4DY6jgYQL3LsqAyy1hQfedwK8
xpem+InNCYCRPqqqXRYN6uZjdRs+B6SbW6B6mWGYzgK/6UCnGrAQp2BqJOp5oqde
J3aD9Ryz7LWZd4DWGVtcwRUWdD2YYibLnNv0iwaOw1RgYI4t+o0hEeoflzl0YAL/
eK/zW5ofnJz9FwoI8SAexmRS1Q0a+LtQPACZwqmkzq7g+Almv9Yy3HDOAsQovNVi
Y7hrY7WdVLfVO6s/qQEUbS8QS6QeoiqtpmUEYHtOu58aUQ1rw4yGt8Q+Dbh++2hr
/5dZTiJUgD7jmKtx2Uu9OVmvDIJklt5s6wRqUwGkRHjCs8SKiGHzxtyH0KrhNy6E
UvbV/KiIuJKPD3sJug1sQh0ABymu8azxHcvJh9Uj2tVGaVI7Aln21I+3t6wR1gUf
AKm6fYlztPQEY4BQDSxrjtGvw1HVfLrUf2/mWgNAK42DOlOm4/RsMy5Vfh1hproj
i2dEa1UlESWCZX3Kfjb4A1Fz7zPe2nsvbaDIaxIBHRP3N4D9aVBSdnKwJ6CEgMkB
m18Mp7Q+Zy+VjAcFh1FVBDgQsKvaM12V/qe6smkvTKRzhT/bVcCQHhhkJtfH49tD
AVL0CfAwiyndHx4fSl6PgNwoz0SFTqq9h1dR+mbOxmhMIDHMoZ9O6xrpLNUa6R8B
WNif5u8yHS7fSnbhoIt0C+/Yn0jdgeVL/cb2o5DMscBsFZQGK9jnaWuYfNyT/WKX
Wdl9BPB9A7QNT+7wjU1GYFlGNACqZmXWZToAz8KmhlhV1aM2duF33/tOC09MbJ7/
Q+FjKdve8nIwYjvuB4dlAEghYcPG9LiFLgAqIDKoSSVlYgZ+VOgH07bpk9aUJvRC
wVYMwP3ZFIqwZBA0EtBOgFvFf37OvGT+1PVS3lO1aaLsxbj7MolcJoVE6nKbJYH3
XBt4fPosoFoen8UFxFSoArm+jNdzMtKPQmpsZ5B7uYn83HZF16zEPOE5IsQxWnqb
0Lz1mx93QDRbH2Utdo72SZeFfGUj8I56oAfo2m29xrg0xfCHmoY4kFx+TznEOQJw
v/Nv0/kIfI/FCrUAsLkeE/GC7L58HKk/OOwyH0BMpwzh213Mdkhrv8GGG1coLYvD
rU09yGO82eqx2YPqB64L0yzXJLsv0r5AMD2ci7ele7F7+BW5xeQP8EY/ixVGU091
ZroacrJ7gDa3Cg2x2lPv7ee3M2pGOuWXMTdXzRtJlQDqT3JJzrutsiFmdxUIf4nm
EcBYyzoZrrXVng7kYUOxMSVPdBkkiC7m6MdRrb9dH0/PUcD3UD3g5hFICTSF6Z/3
FhHgwpVte7xUGQm1+MmDinXTeD06BszLgC2P1hV1f7/JaXFVBc/dBUOUAzLnXLFB
OxAaMx4JMq2DRn4IhMuSU574E5V7g1e7DFgTTSpoebmOJlTUjkw9LlGqrDoLWkaC
b+WoXXRjibLpVg0XotX8+8TXv2aRajvVHWDrTm5lcIzW5tRjPWl+ujYhgIk1Yiwl
p25mTbzLpqxGViX8EWpx238jpL3s2v23toRVrZGlO03vN5adQwarh7NDL+DQyBUr
ZLPcXLVLoShMc2nXsWuGeZlT3aS/oX5iZ17rP4PG+O+h1XOWElHYthXZH47fKu8v
pkAcg4RumlzOkCNMbRvp6Upnd2wWV54YZEAviCqgV/NmPfivg5toScSkqdUoshEy
A3aOLERr0/csvP81Rk0FEEUB8NKpp5GZERnxj5Hqj8NhaeZOZ20gi/wut+TSZxl8
bcL8ZnmWgRgUSOmcKFlAj7vP+cdKWKaGvECoYXKd0L+koZcQVx3o/LF14bkTGJiE
Istuns8w0YQauxfDUFT1kweeako8J3ijf41egLSIJGhUvHqE7EDxrbCQPDDNVa2U
lmYL2OFhPSw8eA7l3gjrX7wSuU96dLL7jFhNjuVxGiu+GH/HgSdal2jr9ykIz5l8
/f6JUTEBJ4CHbW5W/j40+InbdXIDbPBMakl7xwAs19fCmFeBTM2jqBCW8lp9u3gJ
6YacF0UDbNIPQAZwWjT5309nrMHvAroBx/JhtmzPMF8++2Lqk7i3izFakebnMDvy
AQwoi/CfEJtr6wS7wOZOg6gvSJvuxghNe6YYNWupngErsW10XgFr3UMslSyN6Wwa
/OaxPrWG/DR7s/043MVc+KKTz3ySS/CAgvV3izW3afueGWz/+fPyP58Na+/oTsZa
ymfuIpu+cOKmarXHz3aveSsnqJLeJVB7qBqXLce6Leki3S2OJZKAz4rzHZdyLGWx
LRe5F+Kroaltc035lBaa5eZJv5/CbUlRKtrU7JgxrX6bmSs+0M//Da2jp+xE6WIS
fktG6Cpg92lBq4rOvz+wmaB2MRCxgp25FMssQ5Fxqorvga/BzlxivuqTLbHLPF5y
BqCc6iTzD5zCcTZseIz/walcU+RuWk8ASwNkxMgvu4y3L2JMrHVC47gIJaLFg0Qo
vir3budD1kZNtIzCK/O37ENWoU5RcGlopaZz1sx5deoCUB4OonuUACzsNcHGR/GN
n1n7ltnN4fIbYCRwGc6RDzfiDpL5sggHYkt+Z+sqZCZBdS37j7nPfDd0pWb8JgSK
VF8YYrJGSyePdVUuSxzxmzzerQtLcWFIZXPWq1pa8h5t7X7gCzMUbT4ncwLHReNB
p+yKnJiVIS+k34eu3jNo4dTj+JSzNpE00vmdOgjAlOx+71LfNkiM7d7XupnHQtPB
7Xj3c14LQPkBkpdaCoAfWIff6HqaRR7PIRfRM+Sll8rfPyjf1FSxoyIlnX8r7RNJ
1eHbnYyTonNIqo6G476SxLQwKNXHTj9o7e7JpSJuVOlH8TUdqRoZH04BRPL9ZYAJ
mTwPqTpdPVYIar+g5iLdz5YRlw67TFIMRTJ7f3AC2Sesi4+VOZ1r5PJ3u/gNvjIf
Pk/eSLy/Yrz1ZD5WIS4rYCMVAATgnZFKYkAktsWkodHb58DkS+PGrDCtwjLriiMQ
3xXKaelUTFQF7g0fAJ2RqrZiGoy8j6rHs2DgbBTY7gUCtJHa89u8OzIqQLJDZ9mn
YY5uXzn2Pn83Eh7SvqbEBv3m/dwVXeCSe6LfUYeDM5CM9fPFcj7vqUZDEKtOXKjI
gY60zwEGX7Sh1QSNFMhew95LAH6/AjzKIDVQmN43dbEpd79+WS4esGfY+8t/Ym+2
gL8BRZ3ECnyWxxoD6L2KygK7zDZhqCbAvQwtGpbAGe5LNwBZBGSjkDsobToMFhEU
P+TtfyEbsmKlS1EiO5RBM2utTahf3Iylm9UiT5kxBhQmyowfj6VssAKjDbeOUgM7
D+q68f2SS43MDG9pleRyN0/snIQ450EGfeXVeSnGJOBHCWs0x7NxFK+uxkez/aFb
DCKxpvUgCVnoMGl+MuNrad3cfnf4dPb5tQbE0Pl9FtGQDN4vvTEC5fnBA/SW19sh
7OUBI/X94xJDr3O9g06TAjmqtcrT9VWEJbBTg5iCynqRK+bYLajwpEWnaxG9w+IJ
3NpXjfQLSmcS7IcvG/ZfoIjky8FouxvNiK7t+8tqzIiDOHLEaJhSdNGv4ExmQwKX
hePbKPP7HdEyaOEEK0AVGgqROPmlMv9ZX33clRR4TAbkHORxf0xuRcvcM8Ksqw6U
faWGpGuM5ncFPs5oFErg39zJO0uGNvInjqDF/RMhVZkRmX1AP+BWoX60fYisQdZJ
9MzGhUKFdS3qsosyFwu73VitWmcaeo7XY2i86x3ZVxFOY1cIIVkuwVmhHCtbn0cu
B6LYODrwp9mEuHKfk4CAyk3UaYzR5E5x9zDE2NWNeB90ofopg6Dj+rkbl10qOoQh
EWZiHZjbRuAcV0KtJFf6DAhpCB2F8G3rk2YnQCu+TqRyJVYXVk4d3TU5rYxprOzz
E9iNJcXzJcZDG/pvO1raZvbhASDLtMuegj4QmZccBxaX1PQTDcUC9X3fXagf6dqw
b/65zWoiWoPA8eW8LXTi9fGFzLWrbNYBNXe1zsoRf/MN6XATaU0y3YnnvckNKfY5
ztkZBg+G0IvT5IWOQoXXiH0k9uU2jknAEhgWpKhkrzFoHfZVuEXkL7LIK1y67uzt
7NVWT4ibi/fKAEgneoz65BnHFaITpSwH5/0jLA2A2ixpqEwZduuchRulMfeHrYz2
A+65t0PVJOyGkHnx5BW2PSMPdrFNuoC817d3scTcA4Ogn4l1KmATUoWZI9ClHZBF
jJ07ElWSwsmxms3p2h/JJtUW4R9uaUUXgcEBUsRT0ba9Pw2q2prT8ETD2PQlONay
lzPxOQc4kAiF0zsFugGMaK/41nADsnUH8A3djct1grkHiF1QB2gtS16KL8vX57Nw
q3QrzukhX+DsshDHSlpxjL+hANNRwDwwb329gMfcDAk8SFP82MLtWVfHiG5hY5k6
bHH84rF8gk+2r4+5pztCs3x8mys8a1bOWFisIdhTC6N6WKJOiYC90A3jb03RRIuU
2JaLuaMevGX3x34Tm9w/idoXARvKwIeUheMFEgj9bQ5LsjpOfveKUPUOgSQTCJPi
zw8C88U0zP+OI+YLbRtYwsvNTTX5SaFZxnJc5S1v9JM8QwromMgOioicB9g/u7CV
LTTyj4auz3fQo2rjynitO0euF7PZ0haEUKl+NDPZ9BV+9Q+kVGrfaXF1dANCkX+J
kXGaEVNjuTgtL0Aexl5DmOTq0hUtuo6pslZJh80/gs3uuuzgr1JOg1AuXvOuBfVT
y++CJmnUfYXRPLwdZzVeU8Ho6gTgILodDVDeoUStr4mY0jBHBybLuiy64lFvg2J5
Fs600/LERyXswViTF9wOz2YMQDDKSLX4tXFfMMQ6CpXIwxW50/jPnM1Mgx70Cp7p
GTGpqWCpn9vkF7XGRlLmuAO94z9MoGNQB+rHVCFgMZjl0ruImi8up762txs/fsId
MJ5sFq4JKThl5Lv3oSJdIQbMPtefFC0fb4tEX0jf2j6MZEHW0OR6vTyPdcs8TGvU
JHOnPWe9X9h13UUTHut+Bs6bcb+HYFti5aTE5y0JcsBmTX6VHUZ8yj+yxCQyAfiI
itfSSQPfvuEkAxxCmiNKMykvVJY+bJhuu3NQgzWSyDCtzfNCwSn5PVtzcEHf4fw8
cDp9iw8Ikj21Y7B12EL2aqgJNtlPe1XMSwhPqXOEl5ymgonPZyoXs0IN5iUVCRWQ
X7JCuBLIsCUeh01sy0h2gs15WjCDJMiDyZ1nSxCQptODDgF3VCLiloSdUfw6NXvS
qqEGWScRg5+Aw43wHbT0x3I5WkksH5bgS499+Bta+LWvjKKOoxKNXiqBGxwfTsCC
rth+cOsOhDtr3p5hbgVQBdhdIL24Iokej+Bg//aBlJXQmKe0cLaedodka9Ji12iJ
mL4mnquj52M1lwm6R7CT5NDACpkOa39GQdXXa6ebdAMYaw3QgngJoIZJWHZa1IYO
tnozOWhSOMI1aq4Jdn87HjWzDVzeZvDPZxciU1nnqML7rZLeFtvFYx7kZc33Xp6Y
SmwjB1bvMeDVZiTuE8CA/QNkh23GnRDDofOHpNZg/lQ8F735fGhpnHQmiU9Y7sQd
u4OHZy1okFEbK14T4i4nM0E7u45kp2tiO6HgWyqwStxRbSxi7nQY6G3pgrnOo8bi
e5Pp7mRAhsaMjBNAZao/BDZ+0FWMCP3P9zu5N+kn/ALcqJUwkmaEoh4j1nmohkoY
+hsFsjcij3PM874hMkFjfcjf+6AN/Uj8veODbmCKxKXt9RCnPZpjTjRRwM8i6j41
MUvybE8lgRgNHUXYNiEh+IaOpBxKfZaA5DUNYH8MSs3acwsg67qQQeYaJSyEhGZB
SpnQ5lO1TB6KRu7gmj8iqUyDrAiZ23X6x2JHIjeovKD9UABpDN8fTX+efXuVCjLI
InRsJf9v7E2ofMp8agTpD70O7MJS78QqY51gNJFoIjtDmWLEe0g/vPD5T6smw/A2
7UriLdxZekSH5lqVjWnqmEfqUjcYM3CMvPeZpxP0Zwk1z1Ejt4EGPVH0OnfGf0bH
Rds0modhgUtAnAzN3R4IzJiOSoCoeTSL3lhiw6sQTagUzCQ4vjFUQk0GKkd7G/HK
eQoSeDUgrBN0WdO5bvuVB8We6bsRcSZiSEhy2T45W1xPXGs9DmBpn/kgzBy2P4m+
QykQWmGfTK5rP1DnXSxqjNXMf5iHCy34uPDZ8RYu6DpstjT+qysfZ4LFb1oyV6ZT
qEsIsOQbUZ//lo4bWiUQkcPmK8vAXxps6DvnU09DtUR2TxMmLv7SvYWVQWckiFQP
O1vagTXdH1nhXTFn+czqJFz5DNnM1DfeMopZJQQlV47e96mZ8CQIPnnR7BNO3EqT
g17L1MuF8yQYFpn023WJi/crt9uNaJlOUJeKkUO3ZrIJDC0FFuIr+P+nwXmgnKHu
OeySqJhJNCnOX2Ux6k91wsq0Bt0CLykvAqIQXQ82jlCsQQ8cxLIdUNDzyCLcB5pu
ZGZ7vuXHomAPzh5Xbo9gMr4MoEhowcwZRtcJBG3m0OkCr4YgkQlrqLlJUOnE47Lh
/vxyTYI3KvjIfGeQE72VeAJ7t9P8nia8wYQ4I5H8onYp+J6AxBrbPdBSjaKWZEEc
ea7XUov2RQeaL5fBVeoKjS2O+M7Xfw2b29JwH8qyGgWqWirGnk/bnONvu8lESdMi
swVXucA5ocxlGpEfF5w4wKmmCB82YAeeMdyIYIB/MbJDu3dLIbWPOu58wNhB5Uxw
Q0e5KaKAT5k23ODgJHYY07pCpBBue18Vk9RcQV+pOQxRJm0SqTXqKiI1k5OtMTUC
0mwz4PQGg7me3j+J2z3BIcGulNLbzR43l/3AH5f/FldwYHK/8TcteO2PYLawXEdu
ASowEBDMbDaBtx7LFmeJLUBO3X3f8oL/ws6ifNoDmEigYyHfkLdfWEtxhjg9I2B4
k7W+t/2s5LYNeSMXcSyLsSn/e+h74C3Kgrdt1IcTUcQ6uh9cNIo6g3h232ajumty
fwxJmtQVWkI9JgU/0FcxZ5P2r2b16o2PMRe+kHBWoQNbRbyYBvp4gI1BWLEnzxI+
y7Rs4dwm8dC9o4tJlSRNn84iLF8EPA5i0LMG3JczW+M6/XBPiioP0jpMfll0Kd2z
qDAE9rnO6mEq3S7f8QuGF3UNGBQ91IBcSnVQU6w1EAV/G5QblQLPu6UEX9KQfhs5
cWujH/RcL8cg7cx+e7qrPNpiyPT4kRz6s1PLMYy903yCmMIDNZsXhFi3ApTzHghf
rI7haaYLbHkOxf20ED8E0sur+N0HYkKYwJr+v76MaPRMSCf26gyjpiCDEVT2fQhW
8LNstPFHYaKOh/QzzJpYiWD7GSX2t/5DnLfTHUKZw475qTOpN+h5cb7KyV9erJAr
ezpRAUX+Saou+NQBf+tuYyBIqAkAvbpzbwEQCbnpq2Me7xZTbZYMSUN/qU1qHnDA
grmOnzj98FCtmoF1Nc+idTXUJl26fWIAvYdEwjTo4hVuLyYXbF00Zw6vDMQqGruO
1KomRGGcC0oWXxb6mK/Msaj6kQCbmQ7GEdWyy5OG7MWedjd2nxk57CWmBCbTkENf
TF+83M6j8dfFHZcIE669jJUboKuKfrJ+UVYCK+wuXEIJYfM66VIBpfyvRLoB98bJ
do5N1Vw/BsXrRNOxpb1C0YyzwtE+SIRvlCl8HgCg3r1Slpnr79ncX2ofbNiFiFDz
augQEbV9bUak2qeHiNGxI/gC+vJUwOkznaYwMHa1r+QLjj5+TMw01MlGgNSSY/KU
ydp8YS3gOkTzXJYcmpE2gsq2xipKYkz3fqp8WhMAsrlo43ZbbTe9N7/o90ht4w/p
cpfR1ms9Kd5AzTs9IkJICQ9J+Chm0PQIXSfby6LEMs1PZjj1uqA6KBOUyrlHtA0q
x7BRgiS1lzyuUQ8ZugK1VmP4xNvIbkmclXzyZ8T+oRb/qdnI/t5a6eXLXd1ATOc+
cti5jm8zuOVZ+YHglljyqNqNfoI88wsf+ns1LScVBWuIU0L976cQHtfLEX9V7tHU
KQ+DqWzr7u5Kz7fBRYBkA3748CazJU4U0uDA3N2fDUyntq/nvjYvg5m52jDTQNil
uyScIROIpKTrmnQFfL85di2tWKL205h4jC1GB9B2ZQhPbkJRSQLzmMxFsqoQjzhG
b+r8rEIv9Uz5VKcGs/NagSXj4gqCeBUwCVVeZP5Vkpq37Xow2CZ6k8G62+iBiXk4
4+k6xoY7qzM1iGEi5g3KACJm4K+rdyCCOn0z6Tjl/aIDZwYHFjk/M/Zh3KzwQ8a3
6FOcyGlOOf8iHbHH9bFV4Na2qRBJRljDL3msGdLfjWbwPX6RwLBs0CvNm1mYlUnF
FOux8QhWpfuNDP0glqi4myEsKciEkclCM9ODtic1jhPVbjA1w/8E7dFAGAt4uXJ0
6e8mjwkCHDdiGZWjSTChsKoBeiw6H/4BIZib4jIWCkta/7C4KglKA3I98wNS8bew
w93mlDoExYrlrH/F2s96kd8CIGTlRI2UHUt1RvBeLaiiRKzHvlhUYptQNYBuk5Eo
7rjg6EtPjA6K4ZHsqwR79uK8sxpA1roV9DSpCLGnsdL8ufNkU729ih1VwxcGfkU5
pjBRU9vKR3qhadksYwqbLsyXARE9lv0yltRsi85D/IGLtAj7KNa46q/mxUSGBXwS
tQi+oZV6QCMiZc8IZYY6O4la9fxlAz/qL+N91VuU9y7Zt/bXZ+lHwJlpEFbpmkrA
B+S64cqXTqTjDPNiDJ/YVDsbKAMuakY/wBzzWtOIDcTS8DWBUs9hqSNeaASpo/Bg
IJCoDlraa5FtMX9JaYC18KPMxbOg3N0sT1lXPr+Lcz4OgSfJO73JoWmeVtCnO5zB
gRlmiaCblVHy527LvBf0EequCKg8YTzz77UGw0w4CODdlE0F0M6xi9GZabbVg7M7
sjSAH9LQxeRh81k1UI/cbM9iNzdOktyUTByw1WxYmDxITDCezRCf+JFUfKIxBwju
+4hz8VcFsxZGSQ6mNYqusgVpgNH59pPAdGz4MNsz9ueVs472oLLxYdk2bD1b3/1a
1jj/6EBIZO+Il0ZEaJ8UjvAjanL4/0zSR5Og0jNWlnYg6MK2MBQLfZd/cS2xiKj4
TftAD04oBAPje6Txs7DGF7447WA5sFqljSr7JWWsTmUkwASULKvzX8m9y1yD0z0P
QDHHVlXJDeLAku9uYkFV6+DnrjjOesNNU1vyIt+6KNmBD4O+rX82s3n7MkkoAqdc
ETmer9Y6umA4eYDwME09flfBB+GfRp6fmUEWpAwHst+JWw5hixatDaynJaz+cnkE
Ldm/Z8kvjfvyZEN7fnbORsjxpeL6HPsNb+Gjxiyioccb218yOh1gB1AUxAqsHrOR
hZT/lCFQwBpThnfPfU6wYCF9lp8cfoxYX3pvVBHSsjD1BzUJdL7jtiXWJ1mpxm4m
cpZox8yq4EILE9GH3UzWQG0gZszriOay0rQ5sA/tI+1QNjygeQKzMyNUuYFxdBTO
7kCxUurPahJ6pER9W0cctV2qi5kDwefLCICYL2Yp1yhtYk9A4Cc4ZSBmReTGHjM8
kmwBJR01VybOhmgjRhXQUPtFt5Oq3TP9fPWXUxVIf5j3RoLxKxyVzBS+x1ty65+y
7k/g7HFM5GR/JuOBEzgQ2DV/LPeettdrSQpES04MqKzG2VsMgqDCzNXuIl9d2sjp
EueXI8fBZvyA6sgV7sYis4+tywH5qZjI9v9xr5obNdOOxCKBqqj8mgOVTwxgQFf3
IGYLkM2UwudlzOcAvt8nyskoIG1R1lJqHlCcIq8Y+jgMr7ONT9i6ed/R9Cm1+BSQ
E20aLM1ewWhVFjMSfVF4WlekxErkkptXQsSQ1HHRRXulnIvEoAerqzUtyyvY12ch
t54gwDM3lMdyOk1O08Ricjf3rfhK0ajGzYOL2BqskFbGOv9XAWCpRmzcjQ4lxqyC
0Z9+7ahQcTmpm4f3ud+Rl20L8Wca1eIWMPupTJPVjgHLkIV/zwSpkcDIVcVSkjqs
MiAyEiMoPhYp0K2PPHaCTUqRNfed/qZpDjYyrjisUzzYOlqxy65gL7OfAgYpXIVa
bubiFXUkExjCU8jN6d/kH8PlDgyZA50kmTN5rc7L0vcmm2GAhgTT3zWfg00kYb3G
VGXFe8HdLdkIZsMKSsW8OuZZMMuz7fViEZuxfGNxrRtTOU0Wh8HVn8y6gBq3vn74
Eg/MNgRY6cSEncJ/LSU7AlhGzXITHmWItE/kT9Ne2f/AOxfZjd1oMFC8pW81TCCW
m6oa1w2XsA4t4BDnElk76WFTjSVuadnIUEpkR35PWnh22r1f+uRMgqWxWCgGqJM/
rUhUqN7S/QLeJI4J/dBSPpAFd9ogPdjNR5WAVONW08WJDOEdCw8tb4Irx6LLAvn3
+KLJEMlSlQjeqQxzH0cX1Et5yx78WW+xAN8thXZbXllheSbzWLuRuiu82ISGSVoK
APkVn2VuptF3oV0QV77S81l5rW9JRZmnFhDvjhdZC9031harixtQpi0IT5pqKjaK
6b6/fy1KqyhuTHY28tsW9Rm01iSA4D307BoldwZVpTZXKYMw9r3kRQgaYpdsuZ3E
bT+JEaIaMt+ujlIE2BKcNV44GMbbIUrV85nt6yGDDzT/0ZXg+AC9w412mp67zWyx
0ZLGdI08JrYG/qAt63GZraf4J0PYJuZy41F9RToHWO57Y9cJTmA7cE9mz5D4E4d+
k8hSR3D+fXtKYy/D0cQU8ISBy7FdYIpay/iV7i170WhekKbNdOUARcMpgJWu7biY
hlVSGQhMsSwT3tEPiXNKoZa8owCU+Dyp75DIRety8o5UmWwirn7Rr8+ZdXhO2Bvg
qxsT1GfOKamgC/trWVipFJPBYQgRyUyZAzPun87dnGF7ZjaEk/ZR2QzVCo4X1mz/
2Rk07HOojo8WYqy821qM9cEjwpxAGCpZb89Z/WMx7MWlniPdtkwcB+JfCpoDtFvC
N2jcrpgJODI6XhnsVerOceJ87ZXrr7VeRFylAaE++AKRG/lX4dqz2+brBpdG+LSC
dLs+c3tlXlI5tAz33ysti381mE39nWIi2ayc9HbXjQn9XnIif9JUEUlJi1ctZx3Y
01wgMSyfBW5jpnWln7l0bLl/b32rOQbc4gTMItZ8sE2QIapW5HUelzemou4KEUeF
6cj82vsbODzQ5esN5XmupPNp4OJT3xXp0ejlVGZeopbgNlaBiAHGaidiF85uBVee
Z442XehkrPVwnc9uMIQLrPpGYzEPtpK144+n1/XmusxCPPp+oVuLPs/A04uZ+2QQ
WKL21UMoGtIrQCpU5IyAQAUqWUBvEkD2g9Dqvjfp2wPD8gJZ0inV9NOzp3RRC6mb
SkO8OEj1JbRjbr8gR09FAEddA70zfBEgPgMH6p1V8Jit8CAO4SNDo1fNLn9hIdfU
bGma89xI8IX8zKQF038D2yFgqtuCUv7Je4bXPDLpUsobwD+xn0o5BT77A98md1Ha
8jpHp6W6dH7KUP6Gt8dBJezhrtF62AjaRh74E0utRCq79yYZo8VF9FpHs8AjYJnX
2Z0dQxD1hvI7Uh06jrY60R7UZBCgLnAPVqd2eUJCG06uls56uhz3QnL4ZQShZvyJ
L+NXbOAwjScI85oGSZLBDZ0+IaP3BHiHJQ8G3qqJq34UDnFVwAuAiIoCm5KpWuM3
SEeE4uVqGjYx8aTjLozcgERscorkiRmOGNbaWGq9o5IJkp+ZadOEPVXyat3sySpA
pg1j7Wbb9d0uPf0Uq/iTe9O9QYc8eYMrFWDtjwKZgJsRnTsWGEGsd+AnU7V3mEm+
X63meAeUgJjj4rz04LA+GBiQaTPXZByX6UVPDRGmFFHKVtepMls8sIBUR8AQzpPh
cjlnjvOW9+WW+d/OPAuIGfmBBbwVAzIU8+LoBGpWVw/x9fFmmqxo7MeiaPYosEto
69brgqzXJKdmOMEED0phWuKsq1MrJowqL6m9sj5TzIbFvvMs6hOZDuBAwKABhn4a
sotOAVkEBVYruUB6Y/vJQa1VJVQ9UfRaRpMbawsU9cxG6GHCWQB2jPutHU2QIVmS
6yeYMGXiL6nLczUBPh5syXHdJDkUxQrIxUjgGE0RS+Q27xCj+r4a09ak/nk7JmeH
sPjz/gCB4x5Tb4JE4CegBQA2GQbjiK6/YlT+/1A1EqDi2nYWCgvlAjBqz3wghJjD
hDLEzz52eP0XDgGMch3746Sg4ej6uXmOcblZzbsgQaugWHuKIXh/Hjlz8PlnN86L
7nCQ3LJ2zjdNh4yWAf5XpqWpjA0DfPb5MiWz6yjAY+82Dd+8q+kYYscZLqV/zS1m
d30ZlB+95u4MncTl/zhtxMFZtalsS1DZ2MoHtpVeFVXZFyRWQRMq9T8J+1Qm+n12
5kJGl0O9WBaEdXR7LQuZQTC3JgCY2uqlpPbhkmU7bi81asntGwujx/WLJecQazM2
+jraowgkd1DU2dgi3P5MOs46oPZyDUibL5jnB7ZA7nwx176Y6qOhfcR0uYUbVXel
2uY5UKQiE5+O+gEijLqC2FbOkB/jdr6Q9rw/oMbE4YGgRCR5tKZi8/p1xLlIy45Q
OslWY+5yu2dBYVXwIzoaAL8UZ/Q8m+V8duPc9RQMdr/csZ/J5Y7xTCm63zRMc7tc
wZVLXpwFjJWX0Zuo2+/8rJP0abExeiQv2U9ZvWxlxtKF2koW7cqZicdSaamYLdN/
/VT/fMWy24SFpe6F9guoBZNE7xoHFB3b9/x1SF3hwRlWVCEo7MD34QSKD4SF+K8F
OuLDKcRRW+xzeFqPfH+SgmUkoPvImV/xw0CxmtrVbi4cSWhU6qtKRwGJRyw3VC/T
2ZJTziYug2tnrnNxMEyGbqIP7TV12v2wmgp+rm64gPMu8rLHI92TM8e/aJMP+ZaH
S9nSKal/tRVxyS4P7Ny8Fkny1381TzBLXqDgpwbUXY+9vh0EWgCNBIvRpSy5GPKs
ppfW2kqs8KEPtcO6XMp2VcFeBRlQnlyWv3ProyNNl4v9lSywwLG/RoDCCvQWA1XT
Nwfm+fqWLwAOjuZOHfDO3gsGwIkuRpXB6YDf/vqoCeL2Uhqj5nz0KFMzJT+zQJLG
uXTwB7zpGkU7b9GE2dRPW9qJ9Y25WKSS38lY8SYCexHDjPWQeo6jQZG4iVg7Pqmw
0RvTdCQ4AUG9iooVs82w7sWLrXLzq8QGZwy4jZoyKzIfVA37XgTdN9Bdj9QAEKyW
knpqEq07i89Xie89lzJiCDsGAOz5yJuYM//oV15lOsjEffLYZxVouOE48/dq2109
gIxpSb4Ew9hRqhd7kBKxMXG7GblFwzyMzu69m6SGtluEPfwmtFty2XDBm7HLhbl3
c/b4PO9Y8UjPC6vk62vWFIkS5XAd9yIoi4Sp9sMSbJc/T28+/HlehAwZwTuMGrnN
8BnhgtFCdiQ8dxdh+vklO6N+toLA8gmVZWQc75MMhc8ctiNep6w4F6ZQKPimd2SJ
9i38aqUhkqY6r/rqG8XBJRbbeTqTUU/eq9P+4ccmRaIXkoBRFEm52wglWyMjQzmB
KLduy1a3koixPVNQMKnwRa1q2IbK2f0UKBf8HRLRDQXGEaiSo5uxlmZfY5C5H5ge
U48g8jZMmzo0t3ropIQrAXsUf+AQ3LLKJXu0xd4lYk9eO9OzYgsGE7rxliISNxcQ
0e98IO2p1+fh8jqcUSs4uFbMVxB1zGPJxSj0ozN/xllyDzkhWfwb0TTEYOPlLwAC
A8beokqsq0QIH1j4gD9Zd49BjFNpmM209z+p/u2KrhEZKsNrBPXTmQ/1sM/J8SYk
Km9FXLAGuIOl8uMtoubvPTWTZE4t4iVUstznK0tMPAL7IdhnnTCvVhSaC9J6re5L
PrHec2LPLQ9ncZnfcbKLIV52bD4u0YwlzQg8v+1Sgi/8AbLb8NRy9LrWqKLFSolw
Zd0SmpplGqhRYbn2iibJ9Sc+mFx/YYlVDHQikIgCuaIxZhhzH6cUgKk/q/GnFTj6
2dLXDOaB7qh8oQgVQGKq1S7BghueG3J54MPVvir+a60WQJvDj4XYqnKQY1Ajglhh
TEfYUGwPY1wlG8/S8Bw4zWwTS8vZ5iG+3y4sZrFl4AQqp5unfSldFX1gELDM0gY7
bY+qEnkYcfKCnFpeas/9uXaGgRWQ5fubQjGqx3VErIKl806SidE2y7G2Nyp/qiOw
PyV3EbEzYI/ak6BHzwDfqaSv58rbyoHjVZuQjS75KP6Aa5L90ofvhJ3xhUZ5+r7c
Oy8J1LWMiyTXZUqMspt0D6xZTIP4/Qnrg9PrWbpDPQi4iy9viNfTesBIYY9FFRb+
SwDW1LCFog+FPmupZ4r4uLYJRAopN5zmUIqgM+W4hhqfSfity/ogzBNUy4fforn0
Idk/87VEpDRe5mmdWoTr5ZPAthVZh5CbaLiyYmb4bnjpzws9jJYIRUDmqwjJPFP9
OlmK2ar0+UpAzfwoFzRrpuSKj0FKZtY9b8f8HlwDRhX7vzTgsSPIP4xOEHdqdAyE
dA7MU/5ZL0cREo/SiX3P24U/D7yFE1PqpK1eplzKAH6vvc5JECEdvu+f6RHaGU9A
c6SW/8Av9tCiYZ3bSC+l1l4spT2XfxLpgx4u+gaX3qwiQi+lPUWaiElG75IuuqsS
GwZ1FKO8DUcxcKhtFQoCZHgI59deiepFcg+1QoXHsC6exF8NiijJVx2CZgCDQ+8I
9tLNLuQ8eJYyPxYFdMl+N3yuVk2voi9SPV7GDezx+qI4UL1F1si19dQMrzNodUyO
ZP9qrwdFBqgqhX9lG6s4fI0SvdISyKBSzlfOiUHdjlzTJ6hsdawKB3HDMk5J74L4
93DlZVRb+mPqKCscZR2ZrAnIepJRK6tiRd4qOiiYwKX/V2NwREU2OhtV+GeKTo7r
ZXPKFc3RyVx0uHERTcBCr132o65Abq0HHKSOL9Nl3hMp+InDnfTgcx3OmaNQrVZD
vb0nc7Qv6Cgvc6BVQ/y5TT2QqvewLrG9YGm0xFchzjxKjm3LNCrQ79QY3YpNWKx+
WBmxlmhddl+Sg+m4kNte1d+6K3t+xdQAVuzsCbwQggRta2TNsdxG5cwQCXRIS7rU
h7a5csPDvAGS0PNX602LLAc+vE4JZ4JN0X0R2NVzk38DLj1TyQzZYjj4nQo/Xvrf
aw8vNz2ckjU4wZYwe79FdoaQaPvfu5j0CPDoly0HkgA9vazJXuRfv+BOOAA9PN/7
Enz2QZd5jwEbGJ4pDaXesX17PrVg0JhxOzOaz3TffKxG2gCiXU++/pjV+a7m2Y7k
oPd8aXp8B3xCQs2b+YHg0E5OsodUbOKU5PQdDwhP30tWWbAeRPLy6PQ8gArdklNe
koGCuxLGeKP8Z/ID4vECSuOgz6ynO0At3vwwxfgLU8yk1nsQ60MlCf2uWliyvFmK
Xios92xuIZ10wcEMqJHL+FWwr+iSFZbfD8QnmLN+pyLghVLlqJWp4RnoeYeaWkUo
e7WyhxF6y0W2i9s2FLh+QXPi9lTUpWyMkX69bFnV1/q/2IOynaEE5pQfPWvan/4Z
YwqnEYfHUKxl7x8wmK5kfbgu1z+aKeZXlRU4Xnr75rtbQLCe5mSQFoL/9cQJnAhZ
FADUUx9s4S/0QCoKX07O1TLQx0KdfE44sAWya1wgZI3hgDcAPCtgWORYwy1GBlQ4
tJNv1XoH9dNAgpvJpGrxVIEu5sXI3EpUAV89QBkZQfmoyZwRd3sx6nE/RUc/hlSQ
DoXIzkEj2T6oN8/DxDy7mYP7Q+47f8RCErzwwhRDFlOoHsHgK6ZFtSodwUXrk+tJ
CCwJSAGJMYunEgxQ628UD81e6PraM50IEIFCgdGhYqxcv8U8p2Q9PwYG1azi90bv
adlCpM0XfRRxtV5/UMFnBadIof7v9RnKysBV36bHwfIqWIwPJVuOlaAISip4vxkn
z1QAfwQs0mtikShaHnz7wNeK5nYc3uIWOBOLvRcM1IxK+1ubBRxeXdurZNhiFEv8
945FrD8x9fkw26+HkDkmg4R2y3q5/Rri6MdewIKFQj2yDDMd76u0rW2efU9uySdc
hfDcbVL4QN2RxST5ZB3PTpLkEndDXptd9zsg8Osqnmt1sHHBIk0opHl5Ee0ZFqbZ
U/wnP5XgQ9h6DeIbzXFTP1OJexpfpooahcqTU0Mt6aLtlKJxtNiNJubdNmH4HlZY
38WhWFPFs7uvciUhoAhD1mkCYMhzZtH2Lts6bK6NLpVjZDC/4jy2KjWzlZdYiARS
3xr2vTroE+8jKUNkbZku8rvRefLSu36PSqNReWa6IY4IKRouAPUK0m5QIvwfRZS4
EGEbTbNS957o1pF2jNGLZuoYgreY7Oh+U5X9Jod/GgLTry4+MHOLagmu0UGXXHp8
AaboIvy4Zu0/2yXMX8fjgiKO70cikL/UCchxVMdj+zb1XrOURd7S3tEBw7TLjdEZ
SjSvNDOVKkkRM10eHaQfhTU68dz8GAL6Eb57e2GRyiAES8e1MP5ReGg3xi2cK4YB
wYxnQlvVXHn7i8E47vQHWsZcPXnS5tdiTeTDyEH5UbPXfbXCNoH1+O+iK2oNzlgh
VnRoF1F7HLc2SOl//meiJC9SbJyHbxARcG5zuNCjuxwUeKRT/EkHXWophA7Zwcue
dfOEmz2fQm/wXSNxag5JP9Tf/PX6M/1auAe5C2XcdiXLq59WI9tzJK9v2qT1vRRt
YTmK0yi9j3LLYi2/ZfKBDrFokhpQ5pYglyyR0LIfZr0gucgrCjTds2/tVzkJyRQM
aNnLw8Fe++D/WBsxcmnpUHaWKuQScdqfPhIN0YrV9yIDghhJYGcf1cO6VcZxHFgx
4fWOizUUfkb038V4GAPYVovG1GoMvrEEx4DF/hccGQPAcBy1KMiJT0XY9eyxg+dC
w1eINzDMsT/eaELU5eQBn5WmyLU/8pVyYYeua0A3tTYCg0W664pe0xAyWwUF7UzJ
7GaXxPuw6oq9GvZFvcBDtuibfAOtNk4QRMuDVyojAiFLfdA6CJYKo7uiYUmU81Gm
RkfJzNp4trYrHWyxdkjFnsY3OERWNHtLxKZ6HT3FM43yXMEHArpPso/hNN5d7BBs
ffxA8PxLBfyVfUIKEf6fT6eGY+p5h9OZP9SIP2lS/+WLocnV4Q5gR4HHmDG+sf4c
G8apQ0heGK8HTXKRRW0I+Jx4etV6AsuvMrf0qZysYxskLnwugggZbaBHrXB5+OBi
lpQElgsI8/K5rOmUfMqF7yPgUFlxYDoaVQU+ZJEUEZkPPRJB+nrLFNOMkMqIMc+w
ZgNELTfAP8QTFdpLuY2P7YCaOiR0gqrAlFwwkHQnhyrDtsUVL3keB+FC1iFn7TIb
tcoZtOyhnPj1UxUKTrKWlxThwYenFMhX6o0kfTF3tw0iUrmIIRBRNPklPdIqllaJ
SoBDYMc6q9j0OV7mYS1Axd8bj3if+54/i+jS13UwlIQBkzO5+92iWlwMWSQhS4eH
0NVClFsCsYwxY2Bz0NvmuWKWbxltlRvQ8bCQlyvv1tBCIy57xuJo84XETAKEVguX
VAyFOQC6CRTNYa8+Jn8L8DG4N/clnDkR5xXpk7+3yEthzVuSAkoUzUtRGl2lfcNH
91UeiRNeMyhyjc/J/Z3PRlOaGqLzZj3d84TjOEYH+yUlq8cvroZu0lewXuoLOcUc
r4+5SLMYaNXTQJZgKaFqbRl88Rm62v3+nX/OBSQGBkjStKub9wW5ICWislagk/MP
twGlHFCLbo6taz2OmZp+WKU1Mx6E4Zg2+AB58pNtqZzsJnmcgHJRczqngbLjsu5F
JEG+ccDs8CmXyDVSItPfB81BFWc36R5pGwkCyS84xw6vPOO5R3+ZF1UKxadyIvB/
DpjiDeRIokzWeuv2lrqe2QFjew2/klCGK36BDK1aS+sKMamsfTYzIB+3O+zcGMb0
4xNMMUdmsXLXiXTe/na4ofNE230oqJUByzZgsQKsnqKj4WVsHtGE+Xh+1d60ScmL
rgQaVjSYZe/mFKFxOjOX2NCYXXPzXNXLgwPySpy0NWHHL3H/+hSzBRVLoiwvT9wp
SyT/B5cIpyJaDB+R71/KeGkgrYuG1C98DI7i+aQ0oJsnigbKof2EFpa5DX/JG5Kn
5QVybHPnui8+QN8Sr98tszd5WCiufRFhAWbjd+sDHbctlCWRbPDvEnGVScE7105A
r8YKZ9XnNBG8uTUgxK8pyIpParbAHImxscTiOKHdufFTJuU5EdBrFXZSu9+pa1Yw
pahLI4KMWj9i33lcXjTkjbN5OCjgtNRUNs8ZRqQzr3gE4rlbI3OlriTR4M4BEKa+
36g4RHZxwQeSFVRTGWafHrjUSzH8BLcM9s8UfUj+KElo3ChwBOeQjl4jlmP8Vp6B
SAWzXuQm/3e+4RRTE03UEzuCo0Xh8gI0ESebVw4WBXB1pu+OBDo3EL4m8n7CmAYv
OmXb33fAM/1Hw04tiM0nhQmsQJnR9R4uXefBswtjUhmXlPEGrtsFZKDaY7b3q/eE
g3hrUuce5FiOxgDXpbIG5hE0DS4YeYuigcoOPqIj/52AbPBNpT38GNElqIsVvU3+
gxxyBOBYRKj2WOrv5hddO3ULQIaCZZPdMzvEVRxYigzCYjWvMU1QiNn4UHpfOOsC
1xldSBBJHut7laVq7xbgeLbEXH3kM6TnFgx/ECyEZUZwq5t/InVMd187+km+jRYe
v1Ef1BjQr0Ru6wNqsydk5G7ZOeA3F/w6RnzhCXwVUFSmhfxrfBpAWKVzV55Jl57I
EGzjKKyKBiLkO3T5nxA8IkxT7izq1Jx8P/xFYWQ+Mhv+zXn49UdRtjZPj5PW2jo6
1QgrRv+K13z4ABvqPG0lys0SzdqyMyDgngbCV81mwSI8TmJpy4ttXH+T20IMuXJb
eW5MG/nqk1o5YjunZTtSaqCrJzP5LR+vnMX78dOWPMwEkfeLYWKkPLVDoDiNrcYA
TNB8sOvKexrMaFOTX/vQfIRnrLNRIEVhnlJbLRhSKI5WULLWSTnvDTONbZSAB90F
NBQDsMSvqTGg7AJKwuBoMJz8dtKDoy12nBN8Eb5qin6MQW3z5zHDCShiIj/p4mdt
o+x3NlxMi1s9cXW2QNo0j+t8UAnFUL5pEDdHAm0n64RtfFkQCDDJaNlEiod0kn/2
kGN703hisPpqFBdIMl8kmZAaAqE1mBvMBdoc9hBcWu7D3HBWHxF4A9tQjcFSSWLZ
0za3yT4BxbxSSxdyiMzQISqorbluFvnk1aau8CXnT5W5ZCj4XbMFHJorDuIHCTWA
g6AF4+VKq0cwj/MoExppR+XM4CzbKzZxZOE9BfAjEfCW5j5/UHKLswljUtMmKLGZ
v88JtCK2aMf6G7pLBrG8w9dnJMOe3cBGKFLJEDaa2+9VVzXv5TZryLeWHUsRs8gz
BNjgpdrOO2Y56FavNWXTebhEtONinZQnTd7b16WdpSMz5lF1xIZI/ZUYWPUOPGuE
5ycbC5bJ8X5D5dy2tPqk7vP9UVSMPWKrgbL6oLtnCdZTpuV45dR7wXjwUciENzpL
VQliadMD/bDJeaT4f8lhH2WY4cAsTaYGnHmzrBVdlVUOhXN8dl/DQrBswOhtzWtL
0mvSa2aZEVf2drH3YfYAExKNAjsoS36/tf8MJ62BHFfoj1OxcYZWmKnLxnQfJZea
NgU2fCqRNjESXBwCkz1e1N6XWDJdq280qi/0RpMxfChdgAJJ2mhW2qQmgRJC/AkF
OgQhGXeLYC55vfanPg+BzEjbhUPIeUUoKtKxKB2xZMyVFOd5Nr78JGHkhy+yUK6u
64AypisN68/OtKFzPcJ8oIbEnz1OmCg9XRKQw9FwLJG8fkTmeXk02R7PyYvMh7eA
AnOfz3Pl5f6GTvwhYCnqkNI6KaqnreYvivClVjyvZDxiPAQFwbIE7VHkBEhb257o
afyhPmfuUBiwoERT9TJae9myf+paOJtQXDeX+coxkhVf7D/zUCbz6L/KDOq1ZSSd
KbWccyCvTYpplQSK2vmVma//RjUylvHpSn3dXTiKR3M0lLEJpUnsrkX8a/aBr5DD
qXtHBfKzAuEuSsGjUqFiWGc8QJDw5zRTAY6agqveq1cQgLeHUVs/q8x3tCNGvLk7
8AIh2HkZCU3KiYIpZWMIbAZ6+OI3f8xkSgNHTH8fjNdi2cqsdcJFFXgBUrh88Wfe
h4tP4icBR1yRnYAd8wNnd6vHeMxrmO/zTiZVfMxlIIbKRW5508TJX3XpayYHDrOF
5OndLL6iy65cDZwzk7qRB0b4OzSjXCDxbwGb9vRF6KtPCINn/Pf1EYFuZAWWWaBO
c7qzHtjhQuP7dHhtPmT6LNtpWXt74JF3MhYElrRhs3mgZgr+qC5mFxitdobq2SHx
mW6jOAR9unkBVwvGPmZuN3qnCWDlyf/CBmW73tNq9vKx11scbHSOGFjqpadPXO2s
bd6+qFrtYjy8lAzPOylP/QYTjlPzt9cJiGvjhXs8SoBo13lszCcaU6Xkz2wB8kwE
D8iav+BpsZxFJqJVls6jGtdL/3anVuFdbBMtd4SU8DFrpPEvBrWlKUJP5Vc/5/IB
s150BE9nXu9Lzw8guBAmagTAfnVu9T0axX+gufqkDlTnUZ8QPIdu7ch156YAR5dM
7rbKLindNnZ2xiIm+SB56Y5EiFtwhfRz9L+gqRYcqajJ838am1qt3bpHWwPO/V/c
bIPocIqHytnWCNLBdX6F1DHAM7A8lEG/JH5bBjoDhR9Ot812Y2Qh8plbrS6Ys1ic
Td+/wicXgUkBa2HQ5C3UlSAE/zygXqfMuJ/Nxl5VOYV+B79Qh15/Vvlh7HSY8SJo
tPEjPMmaLDQLj2RctZ0jUetajQ1/bzQ8/m8r7b5PHS+S/a59sJCwK+O2mXxHd7jX
a3MOw3smg/ycx2Px2ynOnVxLxHPGg4oeOA5kc9b+f1QMhbsOkKA6O1jwF5eerKtC
T2yQhRjZPSLuApq8GGZNR9AqJ9Hm9CW+6rgpLvj0AqBCMPHey4gg0dNvuExxupL2
XAuvMxUP5QLqR4Zt/MAhRfknDjs9rgRzZFHdJ88LogE3my8Cf2/YC5YdEFZesbUM
soT5wfV0bxILotvSAvHRFvPsjdRRkUbnMJwRKFMKvT5qsWO7HKYVICkbJQ2QPfik
CUVaLH7yw11eKv52hmTw5CgZz5UqO6nBhU7qIsZicmvcMNAnToLpPjW1Qnv8oVyb
S0NTlYlXPokYHHATf8jHUycI1JDCxnP1ku17PnnaIneVikCdIPv1F7Fmws/ubi0M
q9pLT28bZGSrJZ0bk842s+qiLuIVZEHRJjiNdzal7L2Bo9KZrCkJtFHC+YsdwwQT
WaSNvuxKXSpKFlsvBJQsqF7rHOZrnSG+95ui07X7cwPAM31ktwQJeIDMc2Z5sd0G
T/17YTK/uvbWbuCKCm2Xg7ZuS1LjDqPUeiM5JHQQfT5tUvLyxnkOzwv2hk5NmBMX
4njLar9baCNSLUPtEhl1GIMfRaMzPmJ91dy03ZKoD4pfwoffDTwqZNm6LngHTJNT
B3tXV4fqGqImeI3L/QGopee37fQ3c4KfrZU7ASVYtJYpu7lRiiz5zpLp80c11KKB
cWRLce4vd4xrr4ZH5LtVYdMXu2RdMp4Vhj4cxO94m8nt5H0eW3x6lqdEzaFZsZpO
ngzqMmt6LWSY4Sj+46LwGmCKYp0KYuGeePRMXCYy/GYirBZzUx7lKP72YvN96eZ2
VJNf/Jw8plEQPM5tvrJC2M7gbLCH9KD4ao5RhuZsv0KzoTozQnrQGFmY3RjtNhtW
bl9W/k9ldt2duddN+LzWBnytC6KOJ3VdSn9XA1uGeLigdjl9axvspqFKMnZ7t5Ef
hbyV5Q0K/Q6WgrZcSmPNG+7PRXBkgRgflwYhI1sB0j4PvuSdl2LPQiFItwgBt8dM
+hshTXPgWZddFHxsC3RLZ2F2pqP1m6LTzLDu/oz3juO/ALI64IFZYTEEg8h4h0De
2dj/qaT2fzG0dzsgi2XW5FOKlVMDd6KdBvbCogTlDJNBozF2ds3BMZBB+s16ALXP
I2atlDNo71s3aW5+oFETa2OwLHl3dkgFJtnLsT/ykoHa03aPUNuJk3YMA0pM4/V7
abkELym5KY6KunhhlbgOYRd1rF9tL3cPMwTds/oJ2hfFxWy+SuHGHvhK9pkouc8a
JACalJQkAcd7EmcUaitzDcuoqz1vrh761+SIwtfQBASboeVl23zqAqA/fFBDJC4d
8HMmdNFkcmT+CVvPn4YyGDT3BG1S89MNd5tN6YVh6P2CZzVaPwSr6b9CM3NvRa3j
hzthyjjVSGDCAtGRiH7XpfK7IitQDBlennPy4+SP1riUSGY51UIMCOjpdOKMNqM9
SPA+OYSD44JA9eJkul+vKMOmpix2/grhEDa/IU9DmUQE93IqXvXkyyf3Np1Wv6vm
xyjWLP9owLqjWvlrYOkt4H3l9jRtIQlLaPxldUPLCpkwMvRQPLN4IdGn1+dXyD4H
T+z/6w6iY+ui4oZD/df4Y9qKZ7MoM9sMRyi6ym4RDeVtsTnZ5Lx7jDCyMNei86/c
h8vXhaDMC5dUH7VZGW3qJ32P0haUM7IYhFM94+XwoFx/3F0YBSVdShdXHTi3raTq
NlzflscfrAonu2HaAUr0JFZgNEdMoLZ/fRccaNqDYuNFa4EQCVK4QHwaEjSuBUOl
mI/rJd8txs6br/7dVKULcO0ix5hn8rucLcy7UhqHsE87dqpVdrNHPS0KPtyF3D3o
3PyjaWUKGV6fhrcwTsONYVsu1bIloeD5ZyBrGeiLeRE52o6DhdqiPXlSYDTgJTNv
zWw/l4WysgP+bu9+pIaYNAfcEKb+YIOu3gHpuX9Yz/f0kgFvb5wClQBXwukl1PqA
94mA8/5zMM3mMaS9YgthK4TqNKwLBHYvsbNFeCspq162USdWQqTnXxMEvV8LQYtO
4Qvasi5yKdJzAcI5LY7Y7WB3PKluE2ixqVGUZre0CtOrWBg37Kh1cyn3+fuiFcBH
seSgzsAH+N6tnFzRlJXZ1DG9IvAG9+S77R85nw88W9BNTnDVU8r15GdoEe3m3DW1
2yFjwAoS4+BmOMmy3nlFt5K8Eb7+0zpChXSe0Nz2C4gOQ+RU6JkUIxadCrVtdyv5
pfjkY5RZ5Kccjq/HUexPZUlbRuMT0s6iVJriEF+NE5CTE/9fRRikS2G019oANSZG
g7/vPdI1gcUCCqb4OZGUa7pJ8/eue8H0a+aTwhVyESY4yCO0p7drkDxgZKrEjI2y
BmDufbA7bg6U4u7Vho6rvPIRGGuBwer7dNa3PMi8XSBlESzk1gQ9vgS+WuxvIEyx
3GULrURXnkA9JNiZHszuTGHmW4SGX4zUi+BnDxpawr55NfdchpjkCSmQAc4S/xiw
hRE81F7Ff1csDy64cUjwjiO18jbPWHEETRcHoHUoZOyA9a1tNVHoqqRfjw6kVcOZ
hMI5VLMHoMPqcwnoDLFySJ7j9E18gF7E5yLZyahEQUnlOd1Gk1tpERtBXaxV5GnS
aXyN3HHTE2bmZzRCijDnO/YpfGsUHqybSoISJgUP6+iJxvINjPGt9D5r6zsLP7Vl
dpRBRcIo2AMiibnqsiVgnRIlc43ivFridlmeckSKuNEXg1Gw475IEb+qKCoeFDSz
Fx8vgAv+cJDeRQh4z5x7gaMgTF17zkUPicGpaZ10uz7DHILdwjL6e6C8Rh/JzRh0
nOrKHYY3bvxHkGn/Wq1Md39sDZVYorKBc2SNwDAYrr7BYXN9IYugyadSAihOIfNF
XtO4nuEWUy1krj/NR5j+p7R0GNXVO2X6lLw9e3fjtk6ErNW+Lw7tgXKraQ02ZhMB
6oOLyYhVDAVu8tQ3hBKYuv6Q4C2K8YJq0GjGndjPYMIXyra6Snm9oxSwh/vkhDTJ
CnLERBCwGOl6hWwTjy8GlCeIW8aS6qDOuzeSyJ0zHxuFJzgnrUBZUAqFS7HoI4T8
cEVyjQnC6GuZAIBOhmKNNsBL0RVVOOwQZl2D60bGaArtgSlR78fxi0B82m4ymCKH
HMpws9CMX5v8fqJrCQFxLZhBTbJX4Mjtv5HJdxc472EdHbMWBZDRWZQe7YJt2IoL
bj0NnSCMWoxFNa2JyHiSESL2JGVZlY5nAD6RslUNJlbL4TX16KKdp11Hn3qiTxhx
uKimWSN4KF1W9koKen8Yf21wIeDzDMNjuo69be+DQRw8/ayuQHr2y+W7npmFbMWC
AepvgANXdAkRVy888IcTbG50dve2V+eZvQAxlg1rcwMl7RspuUYqv9RmshO3KL/r
Ax2r695fS5CvSNPt1aW7k1j37v8CMV/cKYLeJhrdHbPBnICK+RCk3Ucp42unQaEb
jZx2eCqWMqjzREglooIV7t3U+Vk4FEWn/kpC0HRVcY6ZlfrJopCDzL+6p+6g9pMg
a+0e84+zKew/jXPGkENVORHa3AdFIpeOdKbRtfPCHMsPTRNBHeOJ7+50AtGUvPkU
aCvpaxeLRJx/w3cP9jr/6YyVW4Aapx/07Tn3dOx6PhyvUJXF84ovAi21agwPbEQj
oVo24KK+VgujugLqdcm9jiP+npyKoBoczaHt54RLB7BZL4fRr06xTuk/hfIorpBc
kNAQUnSnz+g+Sk33npW6Bg+udaWjwb7qhmwkdHWJD4eQ9FqKLrHBM1uBoT7El14w
9i4kwwrDB0UjJ4k/sT+3agssVu5+fNESmrz3rQ7DP7oAhm1jYKqZDIQWl5H06tG3
NeUUVpfSDFymICyzxsqw7cfw2qYpp5HC2vm71oMd9qrULTPepX4UMY+SJuB00JRC
E0h91TbQSYcB8kXp29KcVLj4un1LO3h/cKzNo/nlXmSWq99n1JY50drinEor0HTd
ctuU8qILOhA9VlEzLxWnbrvEkYEXTEvkC0LlC+vgJWTuOnSC6vtnFmo2JnGQpNmx
aasiAXRYRoX7Y5/UnohEARoNzAkkHm7fmKcQzZ6ydv6bR5eoa22a0yGl0rVhjtft
6/2lU7OVQRWSybva42uGyCzXauJggK5q44IS358y4s1JsJpTA+iCP19D1Io/5CoI
EMgRVoRkzZU8hLMqe/6GJTunL8JcPeWA5POsWxPCovObA7eQUTsI+3o7DFsZHPcW
ZKZiRFwtKZSh5PSWVbZcDZNeijNu8p6zJQhkn7Di4fJEdRAj04Efkd16wZ10uvnR
vQRKXurRcTN3xm4eD2q/8RYMR1tUGCznPKQ8wXwqKs2kLMst+v0TOl/2svjXcQMn
Dz+sBSBqjifJkLW6qUGU+J/FhF4+Y8gjEuUhGYkmUMmI/3G01QWpFokhIoRCUxPA
MgYF1iFhAE6SU6fR592aa68MMDMaU40+A8AYARfa22yWVYzdS/TxYWc9jwGosN03
sEXoyayiatT2Qr9bDM3FBzvl7Wyuv2zIrNdNUNNgQEuD2x17CPtMA6dRZl2TeMsy
dqzcCG5/oX7ta54kxJB/MC0UXV1OBRAWiW4vINFq1SftRph41LXL5I5prBD8IMV0
KtBAQ+IdQLoc/IPsy6N4t33GiSOfbmroAJ+nbOCF/1OiR7m2P/qEej5R2h8Bet3N
blMMh1D1w+RI8dkrfm3kOB5qIZiLBjHGCbiWDnQk8n+fBVmM6cWHKWSt8OLB1rlT
VOo+x/uY6eEVTt4GjEKdvsE2+OJVHc7Qv0IhVkwOykAqc6aYoyJ35nD4iGds1mlQ
Qfqfk8BkuczVDfMHe8gQnNZsWzwoW3SP0Do8QpWGf5hw91hMKg0sHKjIBBkNZp7/
9XQIjRyPAJmDagmwvXAr2vTQZ4sI1v4P4KxTcOzuFRbrTYyWWXiQQCW9bJtnR6s6
N7YtWeO0dtYLnFXQ7RH2E2boe/TylfxijEPi1tqvibp6AqavaziYDCbMxPEaOyV6
BqvQuCce+RmWmrxcboNZHhJWceYsJTl3gbmDCBnLBGd1E6HRFcZqiuEGIWZS2gjE
13HeYG2x+8iylyhrNV/QjhskaTrti5aGSZ5uoeriKS+XCmzU3T316LuStrNVZ1Ik
GyLWGdCSttLfp4/MTmacIszbzsbnw1k0DsNPmzoBZS9H/BTY5d3XF20Rbn/B0F0P
/8pZ4ceGTzs5Uvv2lnZSXExUnOO0EWnaUeMlebGoF5BX6/dVLHBsmtk5L4H/GriY
QyHJTIRgip3WL0S33pdd8vz9pA693NQaVpM+cs71QZZJGpVf5HwAwLJO5SiqbzOw
vuZ+reJprT+qOzb87E9BO/G9LImskeB/VeUHa7QRqICph997AYSvPO2Xo91mj02z
FonQv9o+tRM4WIRaEsGttCQI9bRVCxUqLb4CnXiaijg1qDKkySvAvrBkguH7I1hl
YvpmGN6FZrUOwS6LhNEZj7z7WhB6kIv0VFdPizzxw8uJbGWO61sMI9ESGCOvvgSl
oQL+Hrk8fwOsm4eLVll84dwVBo5dNhxicNILLH52tjMkYs+nCCpuYEm9Ty+ehh6O
CH0ewpQsTVxjW/3XJNyWECjExago51WlF0LXp+43/WHMQsdAyEByeydyEAeJCAN4
FboSrUIruZCWk7JF/QuCYO5B9jA/D9Wj/pFmyRRQznZU0ur5jSxf/aE1TRSVGI6o
qn7VycsDYzL+4V628NgqLCce/Jxms4XK/4jA7xZ93wPql8RKas8/3hQw4lnvGuGk
3cGEonVoEbAdKmZpx2vF8LQvye+3ddd+7IP8jC84fsE+MsQDS6D4r7jNGaALToHb
xcxRRwSMH9GSIu+gQkAAp+tMI3TKZ24kkcf0fVm9OeuOJQUNN3n9hmnqooJfA0VQ
hvDXqi80j9a4m5B4Gv3CNFXpgOchutlFT0oACqR1jDtNfZWmLDj2tXkhvWSUyFoQ
aGmmKx9y1CNEcqpXXLDLW4W4aKoAWdMx0MJ6h70jI7IUdlMXslPddfV3e75ncXoJ
W3+VSFW1Jc0lWLaPyznqnRtdhq6WILoemO8Rvm7Kl1l2D7JcrkT0/P7rY2hJT26v
x0WiDxntk4O+46nLabUQ1dY+Ry5FHCluORDtCqqD1uekkhEi0sqEp1IL4TY/DLm/
fdQoEUKuXCS/vP4sV3fvHpDECFSKoaff+PgeWXr8c3fN2k7LYqR8u2k/LmL0y6J3
RS3yudOsRpjtBTvcUV8kgV3h5lyefZj7VyGfOQTa2s4AM675STsm8EQ4biGv7BR5
4Qhdpkso68iGbCuQ4nFRlCcXSoNCoP7CDkNpLoQX+eqQHgwuKWaZDjc6g6Y7k6y3
JaaT3DI02cdbXklM0a+s/sNBKEe1XCUHMAgSumKvNPJx5dCKuw9/jphTN+SKaqEO
cs0zfG2aQfdhbpVLQeHeVqwkDui+JtMf1UBUrI8WtOKqLTVlnrI6tC8dsJO3oS5+
2XVAlHuZV1b/uWjBKTAcMjwNYquvvfjn1/xxuwb6/2Xuj4dXmyMFhaazJ0pIouUQ
OXu52AlqqLrNW3jKgaPOSSWQEY4zRMSFvDx3yQ5OedfgvVNZYi+USW+OObJI2zqe
rQcpe+4O7cOnJkW8bEZyPcBTQOvWGNbMetLpEUCIMU4ccPUqJRZVArXBepZZz48h
6GSWOge9PzOkIvSRCy+o0NmlPT9I0OCDwT4nIicJz5xvr11BoqXxUSvwyEJOzXGT
4wvjTsWn1SItdZqwrwXjFSBhAt/92sKlMepkaUQY0UdDzuLH9YxCQcosAylSjylN
HuIegyuGpeFEiTQtrcxtHVtNkOR7cAGqlzyyMKNrUz0SuREKkXeJPNJOwYYjPAfk
J+wJypQ3G2BtHXy8vFuJkuOJdHfzfN4o2/B1Q7fHiE7t2GAqqaJXcCv0k8tfu54Q
E43wXULrDAhoXj86Ypx8bU0FWffla/Iq+SU9FtE5Uj6dXMcHzHTUBRt6xG/xQVCU
JaPJd8x9EU8ABP/TOMvE7kZGYm4K0dDHxOXW5/WqpJ7FohDDsNB1lBsGKpwt6FdT
dpFthW5dab4X4OJBWQP1wW21j+4C8u146CPhxSoQxEaPZG7oYFET4uUy1Xm5PQ3A
2hQszEaRW54gmAj2IEvejhm3RbVLu0iUreivW3MNuCpFIA0dTz6835C88sPVz4dK
5ALZdxeMYgBZwKbhmMZvhQhfTl3VESGyJAsx/yPj8B4mlcpniE1mZirh1FS1czlH
mRepSZBZJs82PY6ym3iMX5NJmUFwTCxsCvmlRyDVjUm5DmhRE/1wH1EweharaSLp
24CLUh+4ddFdBKfxAXcUK+JYPp+sBM1Gxv3XFp06eI/Z1eLbnqozrmOtNHPGtdGT
pJC4fgXstlDnfr90oRUrG1XaEHRWpgX/07Tag7BqZy8OFtw+NN/jYSUBAHr5/kcw
sWpNR+q2Zq/9FBm/Xk4tqVDCBqa7Z5Fy646aTkFDY9+lbHZh8uFILtp1X7oBPTy9
EsFpdiHFSg/hD9nFrLB4v3QhK2aA/Q6XJHiM6fRzhZKijiDZyUoi2U4LZhCguKCV
Kbi+guR5WDVWiENtfzLWdtefL/er35UopQcJ4/qz0ptSo5tmJy+QArlx0rBbt7wq
s1mPay0npQLxaGtczL6ENt1jC600KQR47j6mw1I3/h8G/e+Ek9lJefn+9W3iiG4l
jVre1wOEjKNqZVuVXQzyWwamqDSsLqyhhE5zzS8op43ClOtXRCC6HRN4mIF/o9+r
lrO5F0zkmfupYpG7T9Ai9cruFl+Ax0N5h4p36nB0k3Kd0nWPHvfi8jPtrAMl70gC
GGWe66cHdWD4pa7QnI20KbT4F3f6PEuma5W19/5G/uAs/TbQfPkLmJqrtNNS8lo0
U/oxZlXabTMlFeTXQIKp+4zl81We/NUYJWSPACygr7sjB4O75gGveZGcKVMdeGZp
hxMQf+j5I+oIQR5OmVGo4+TT50woMJ1UByFnwxycHSifXJ0cn4Pc57o8N3hvVyxb
sfL4M9za5UQ8s63y97zA7n9Tb+iyfGqnpPWP4GRvy19VdHJhgHiVzLuMQBPZk+65
ftgu9MecK1Ha37L7RWo5BjtqDHEG+XTbxJy1hHp1hIG2vZqhvPfoz6Vw7V36BfGM
1VtBLXPMSeYFbyoVYIM3oqcckh9vHSc4S0q/G+AHYY6rwRjX0GQhur23YLB+F25H
6QxBZA98s0VlHgVSGNB73QLtpWQMamkQ8i2wZM1/FtXD5cCTFixqgmjyPVSRftdI
J51kK9DHjutyBtxGJOuolm5cPUdEN/gyOFkQMFx+1p7VtZSUO8kwjAxcjLA7ZnXU
w9q6Y2NLNfEGEEDa02TmJ2EbZZhTI8gvMXgVHhDJH7JebTIscVbifTL/5J4gfZ5C
23+5UaZptQPosCFm7kMoQ5XKoWVQTlZsg8X/zg7mtwdtrcQTTACWCJLTl2on2z6F
5QDNJtXAwmvOcQLvZoqDzD+gDuajz0G33mwNqkTmUCQZVZnmTrTBU3zTdW4xdewI
HnLrdMI1vIchXIBlaZzw+BeRXzfEpJ4CxXQpPjzIwKoYDUNenIuVCAcSzWYrwjeF
iJK+3jHeCIGXBL5NZimpmZjIeuGGGMpujtsMkJ96avZ0BB+OnKa/8YDAdhdazP/4
bn6aTPk4J0KeRyR++8YMtuiFXVlHpC5GLMJjCS/XN5f0jxEhijBLl5uPD9YsJmum
ZANhHNo0G2hy6U7wqNCbBOH3YoSEWtwoX3gJaC9WXocPT/U9HbQMqTzG0IkeNUp7
ec29BgikbniO6DV+6hoUE3ue9969EG/W4zUYmxLlt/ipJOzirTOTKIC/U1RDdCjt
393seoPzfiRLYevXxtVyOasESKdTD7pDlcbcSWpcHtUptnvmSKj2acWJTAhDD75/
r8Qwk8AO1IRP+JMJ/du+I+5V3e6qb1wfYSkulEAQWuM0xu7L9SH66AKqts6PUdV3
gzqUGM5pHvpNDOg4rWqC1ZxysNCcD9m6flDTDGb/cIEstIHbmVzLAmSr+81QbV5h
SA0wZ9BjgtzdE67tdHnIBnZgqNQ26lnDSX/t2ogQRDxqWIN3zmtFmLPC/VEUCCwM
wUfDtMnOjZ/R+x/ay914apLz7vlUQ7hRJVlPrOza9bDbspd+NbKnz7pMIWcCfOMj
KPQgiVze2MsF8AcotyhCQY63J/GFBVPtrkXnWpKo+og9O727qxF0gCNSG46vD45+
kuwOxzGDNmp94eDJY0ulfkfatDRkW3AoqtXMC04m/tplOqfwCnj+GaC/IitBV9X3
0YIs5Wi3+32EkDBqepV+inlrm9FLFDAveaom8ENM7SJ5hps9pNbsCrK1MVIwdDpJ
a00NOH18rnK+BQ2heUF814R/vJusPxTte6I03twfRuYSEAGEymuyfuYZ/jdZr+ry
J/JLZPxY63CZHG0U0fFxNpqzFglAr6ttuvq92fRTebqnxFNLpRF99EfaoocJZVUA
85NqARRs9vpyn2WtR5TRvfHnZlqkXs9WL3ep3mFcssIKXkdTKssWBTqNfBznaGWC
xanxd0uPIuttJf1rp8fkSFsEEkIJIbI4T62QdJYqXtLvEcH+w6ovpqc8n/Cu2wiY
cKQ4plAeW41Wpgay9degZXPyANz+Pbtk3ceNhXbaRC0KHR8CVaCJ9SqqD4HiRVlu
fif9K6m+RSaN6tzz9+1WhbqQrl0JQc7owAFLAtSG6uS+kSYE+9AErVq1cfuSOOXL
mLIBo+iR6swcVMf0K3Rb9aJjMsSo3NNudIdcuu8td0tFhFWiayTVG67tu2U1IB7o
GtS9VJdj2iUJUOEzo9btp4Qul9hefziZD1phsvIN8Zz5/TivwfEs10i/GJYYcHu2
M52VsGTbhKtPeURbj34xPEkDJbMSekXM/BrwVmuWaSYdAiJJ8q8xFszMDVkSKrlH
b6+wToFVBBQh9K993Xfo42sBPeiE438gTIuoPlqMnNm9gKhV6H1q1WsZsLPug4pQ
PbkZP37KL9LwYf8taypeITGEHYPSMgnd9JxbgT9tixxLN2Q/f004avmPT2/1I9cr
f9GpmIW/XdXShoufBArpTKQnaS3udzUdc0OSsduesEBBx5w7THnaqNqHazvdM0bX
rIVsNy1XbyO9e2sES97dA22Z+PxgalQYcdwu+JhCeFkXf6D5oiR4jzSlRN+UAumP
gisSrPAnDgrOlCVwANl6HUIxs7LR2y5s6vKOz6YPvXf0T0wzeexrisO9aRL8jjbb
yNURl03FrVnn6aE0TZI6Jivkd0e7Dw4wPLXBo6AzQa3PVyaNscxWiNy+LYCOASYQ
9scDVfAdKUx8pQrEuioCY7cQkcv/sEoh1yNlYzn3g/g2OeQvUqKXn/1q/57He2Cy
Em/LKD3CdNOsxgTE5dwNN0GN1wswIhDommB56s95adO4w4bBkwc7YP4Vd7cr9KK8
WjXb6FqkhVUG2pd8xBliGeP5aBagZeHN96SboSh/LIrr/zvVUDKX2sDfPuLjkDI6
AbdLw7uUKqnWeEMhiS8mpRkPsNyOfzJvTYvWR9Ue3/Vw85zHooJA0RxZpndoh/9R
ROp1TpysBXelQ+Xul/Lcpxdo31mt4w3SD8Ft6AgoEFCpUGHVrRoT4RL6oRcn0+uv
0Ht4VIH/ivQ7g5jzIqIr0p6jXcTG0caBTvB0A6FK9Ku87t7aYxAD/fw+zPBfkTSJ
xJHaGIpMyoGXniVqiPWTMrdC09zgwKX1pmaFi14kWFC1TZ4PM/B5NsLloQ3iQbuW
8kWoZOy6KYlgwSe8Es6TI5X0xgaGIgLWU2QG0vtpgeKyW0nyCSJTIxGRPTRrsksj
VbkC28HsHvuiPIPdLkddd90W/XVOBOm9pn/b+Iv+WKApc2W4qw8bJvFd4gCfqpK6
2f/34vuPnWGUvp3w7m88aDn0rHxKrbIBGCG8KT/UCOkwi/yoYvkxCOyAoDfBi4iD
u6n4PFtjD2VPxKZnhJtQnKbr7JsqLAgSXIFwGQWumlbYxWoQyYBb7H4GI6ksDIMV
7yIRzmGdMJe8qXVTl8Sdn0OBWAYbAeUlGngbI+o4qEGjTTQRQ9o9mMBwJJ8mIorT
SwzmS9aDt8oFTv2St8MChvmj/oN5cTIvNtEAsiSYvj1kdDTexSSfD/6WdOKVpnkz
uEPezlB0GBYBM4xyQbdopTSB1xWYOSGMKhhrNOZlhcqANEBK6PVne0/zmiSP4Gyt
AU+nea/xKe1+pxPpw5kVor7/eEA5pwUbkCVyZgX7/g83qpyVVM/Fq6wQ/6tivVE9
sJgEWfAbKCr/hy4H+loHJDtp6q6e3duPPB9oWM1cPJFwdqLeAhDWZdrbnXJVJa6Q
5kouxdl/gkzrqY3T0x2Xlg9j809eksdK7JAz+miGHequ71HhtmNbjQotWXfKFBhQ
wKQY9hWUaEKDMrn75BYzenujE3KG5w6b+234YX9FSKC/xBw67u4paFwIfuwcgUGO
daJQDnBgR/mGJjHGYtIjcb/2fwkjqVY9sp1MkwTkFzdy/0SrzP9a9dwWV3cU/YYY
Tg7Jiu3ogIpRJzAjhyH03DTrf0mLxOw1NrM+C53rbp1Njt8ZddVHK8oPKU93y+3J
+coKgJzWtWOE0+Uqk1UHA0mf5g1XMWNGdbPtfa2xOdatzaO0YdBcKXaCAHHvciQc
zY/jX3VCB63fHjLGiGnhbvFEyD7q3lPiYcDECvH1ysDpei6NeotSGU118HISEOsN
NL7JNew9fOA4FBF4j9SDTc3fjUvrdCb7Js+fe7HnbYUwCMLkddN0mltWBwNKZ6+R
csxtHEhOr813MQC+b82CCeY3h+iOrrtieC3C/xgSO2Jny93DzBE88EzE4i2gcDTa
jgeRO0RBnHIxplavsH42npxZo2dptRcfveUvj0Wc9HCLvQapUeBPR9AewLdKcpKP
4S3kmkDW3533Xo+LOsub3RGs6p5wLJIFGR0607PcVo+IE1xoXitTu/wPpFzdEWJ9
HTdVd8dkZ1R6AgnhHKHx1DML3fNnxsTpXN3ZHxT8FizD7xcWztDx/6Eh1G/Celod
WOGzyzO+6Vbye6wKz68BqiKO0AiWJE3H24zkSjNa7UsN005pP4ogwK6YHfnT1xVJ
YbZIrjCKFjo6UgNvaPN5BUEPJ4FW7LjuW3mLovvqMupV5a8OpE7KeKsiFpA+yqwg
6P6/ujIcZDMVnHp3zaZVDztO4YZL3gLBPEVlzl547xgKKKDOEI7VidGktrfOqx9n
ikbY3Ly//O/ZVgkPEjRqogaOV6dqcwH0y2fyHakeefGIAb5+Xm4Xn/s9gMeZp6cB
FD7ag8nWjr8CYJNTurcD1cIGIwC7tvNha6qZU4Hf21xRk3kLo1ybLziPk0zBAHoc
F84kKFpW+6cXf9Qmg8G7ASaAIAapArBiUvE3Wo9yL9cVLNXcqhfVv+LxIARM+Dyz
ZlgvCrWKhRu4+0e7aROQ/m8T8VLyv8dTbbBw13sNIT/UBtpK7j0aLpZjMWAzXafD
4O+iVheZzCQ4QuSrpHvruQL/4E4El9D3DQa7A5147scaKBu6x9MaXBakhIbpcT90
`pragma protect end_protected

`endif // `ifndef _VF_AXI_XACT_SV_


