//----------------------------------------------------------------------
/**
 * @file vf_axi_hndlr.sv
 * @brief Defines VF AXI interface handler base class.
 */
/*
 * Copyright (C) 2007-2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_HNDLR_SV_
`define _VF_AXI_HNDLR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
BJoPQDUdSvg1UaPhW3S3yxv37XONpwXyAn5KCmfBWLHPs727XcjnV4mM2iaylhH5
kYJucGHj1/liBbfGfu1TZXRSgawmCe4JRAknoTu6AapipaT5lYhInmPXLFkE2Q85
G0dsG92RdYm/GavibXNdVBk5tGRb+611JZ2c7zQekmJO2V/40Yg0TBgR7Vzc/p40
vLuQurpfpywNN15i8ZOcRnqsWszwVLPOGNVwYnsEqf3c0C5c3aAUzTGbIvS4IaV+
/hHvxVyouGHIH2SGhW+b1HHMy9MnnL4UqeAvYT2GUkutZWi+Fxu6350Nc1dYE1bS
ZhvunqOxgBGOaaVaVTYw4w==
`pragma protect data_block
z3xVRvt205zHnRZKk21AeIN7f61YurtqofQXeYndP68v77pJ2mWE44osSmyaJocM
2d7TZNfXAFdaTZLyhCKmV0LkUJmqFkmK57/M2ED5xads5Z/0yYrbN8uIubLZFnwn
o0Gind69S4rYKly/6Z9vHi4gb1X7O/tbpZ/wCuL7m7cxlps3SmYwtFg1hkVXfM86
1eqtYzUxRQioFeUVrzCEcFVG5ZRdMttZOMOJEzqcRTuROlX3VS0x4CPaHkCFNGjd
5fSxtD5S3GN4DFNimiQt04667VtKlagqiy+UWkayQWyhQipY3znpY19HYzo1CVQL
vDmZYYrMWbXQyhpM4XM/JXW1qfEPRc9z+9jxDFWI4cpi1rqQBm50fo8xWo6IvRot
wByTXTemzSBgurgqXbwwXUVm7y3B1OOWV4yPrseKPrU7QHMOUw2QGGMfhtcv6jra
j/I6iY2fHG844CE5vL7bj+M0nQvZLxwIOA4CKWT5aSBiWjb9WemkslM5Awi7ggbf
AI2tto8Qjv2Y8Vt3Ihl5KQG5hWT1tgvxcrbfvYyQTdkNzxm0NGApqo6TVqV33y+c
xLQugOH9yzpkHwWshVDIji886Iu44jAlkkPc0XVVNEmNaPIr069huZOXd4oGk6go
n3jJPE5IWkskomoNs1XrIvucmMuyYMJpYT/wCCRBG4xXxN8zBktHBHypKuVgbOP8
aK09vs5SF/vZ5ma5TxoWQM9G4AVm4b20mnyBZAOGjD/kZvn75Tg36go/nies/rcp
7oZutecZ9VhWYWWcKw1IFNGZNzjgwYEgKOJxrcqo+ac9VVzp6vKeMm7eFmbK4aK9
4/qhYeSULQSq8sy2PDRErQDHiJ79hgMg/kyhiAbXG//x42IUODwskYVRcwNpe2SY
KG9r4t/2ejNk37JnNuAkZobBVisXlIVPUVmomgyRrKWR/6Lhrn/pnWEPkN3BLVk4
R5GI7yTI4Dw/NoOxq7dgCMYrwy20yoRkU0cBvWCx2kWw9SLrBS1EiJOODFFUjz5c
7otz/NVXQBfJR4uYPPCM6HCxi5GZFqWkfx5opSfvop98nIjVAzc1RQxkruPD9eTv
v8weTjci3VgS8uoTvTecqAweUHiX8rAgRS8Re05OIl8ro+BIoMRVTuNI/zO+FsuW
Azv9WhKv1W/4Y0Z0lh/JJTBtHdsr2Me2iqdQ/nJgQd4u7LZ+pQFmfuOe4bwyTnkx
CEyimEl1hQUx/OZ5wDAVeNULudhzrp1gjiigc4EkuQN1CtxWzoY586N2ByH1aOF8
CTESyFDz0E/8+Znx+v5k6+3uYnBxjKgyuJrzMyXVO6+yY98JUdURu9aKgoOmzxda
Myh6MaU1Yr2RWsDQ3KCC2UDaCEkWLeLTHyg7Njf+gcsUYd7AsCTlHinoizQLKuY9
xQWQnldEalPY12Zpv3UENqN4sI5N05WvbOMQyjUc1AkdW4dO+1gcRIob+kU4/F0V
nJ7WEqM6+jP7VeZ8Acdoli2F1vZrqWgOKp1gOm9gduMikmjqwmbdfINuC3g5ylR3
VcKTRIAH5RCtSerlJl9ASvQKpf4ITJhSdpXMtr++AJYi13R3TL/0zCkzKre+or2I
SLWXForLDqqy+VoB+BfZgBxxhG62rgYDOHv76oXBKfy5O9qgpOM2dUIjaC/1LCj+
O5MTC75MSMSthkOqB99csFxxjtCtD5EVO4A12bKOFu/+Axh9nne4u12SOyW4XS5p
7L/LJ16VJl0S7j+jzNrXA/fMycRDYIJ/WTqBJCs6k6iJxP5u0alGy6gxKIQWjDoF
Tx0rJRrBZxDHf1vkyBIoYCZaMU2ttycWSKFneWyxK0xXAvh3JGjRI4g0o6O9UReQ
vNn3o3uHqcJ/JWExSWbTGjr1Rfi/sJVPN5hSM6TaIa8EGzj9t7ytI3fNsKm5VVNV
jAxQA1b1xKxRtpj6veLf9Mm8Fi++VQwCCRvsJaIobTgBSXhgITYS+iAoKHmTlh/L
Uqu7VnceR7+SBNIxHdAhFu1t0jb8YWJzX3/5ouV5LsIb2FxXBfmb+e3Q4OiSMmpl
1r3pr3cbJczmNiWFHiL0NCbZ3MWM0jUzMLu3m0FbPAIIMN8VV2jnYK48lE8GabRC
IJ72FheH49sS0cFQLB6205WHC3igYQwEcy/GxlHJpQAA6u/aPow2/Kx269erJDue
DVLYMCJ7jN5eZesMEbc1evToUA+q22bQHhl0pn0afERjqxWVeLj0Qi1OHjYrHBK9
irqGDexMMw67aova27oDS0dPtwJCiwFJMg8uH8Ws2msH4p3VrqrXmpqH0tWSRMMp
KUUhX+oi+1VVXgTv0oTImBQVAKiUMUX2lytChukqPRmhA4ra7ky1KkSr320wUYAi
fJtMtdqchVnrc8sFIG+pQ+nVnLiRD8yV/zNo4vVgDTQ0jHcFa//fDAdXjyoIVfxh
28Om6tO65gZHCj7A7kDQBqEkDqrAckOIv/hwNlUZyFIf2BpAbCInfyFdGWkyvjNG
ZODb32DIVrR4bfiw0vLDAzwAT53giYVLSUBBaiO0nxuvE4xNtPcrSTdSMZFqCuH9
qaa6xctm9DHEwmyzYJ3jOIClv+dJ4YS2Q+8SXtboDt6PKc+tdVkPsGAZbHX5O6zU
hDarSPMoQ5kFt6Rlr17jmLdbVAkE6M+5yAc/FrGEXBly26mAis9Xj6DeaVqs0a6d
GWp3qRsf3sQfhYjRxTYOSZoYA66F4Urv3OSf2Dr1kcpBbRIY36XnvenMWU6Q4mGG
t1l+2mUHmnIBiVDfBd5/CpDq2WMR9eYdeylBLUllQRVldiWFpemwDdFvtb3B0QRl
Z/dyzB5quBy7NMOhdEqZthmncRR+q/kv/ir6seJSs26Q2TWbpmduUCjjZnbk1JgA
XC8TXgT8wYwBXnIk44kV8ceYJbQ5qXlxgaT+s4iZf8PrKxOReMs27WNxZA1I7gGs
PV/sLK27isprcLpUdZiOhWVj1riYXJeI2u0vDj+p0ePi2cjZ2JEJIsikpa7CBA+G
lwW0DbyPrr1imKU1FZZ0mhv3/FZxp9PoNnbju/WKv+77tX/nK5htJPVhKfpfhT8o
ijWijHVNNSR5tsLAspQr9SfiJ+pRCk0bk2oPv9TYuj2wBGigyhWxo1xHShMVwmWp
mqoRBe8G3WViM60Gm1njOravLtZQLkaNgEUFo+MVwLMP91X6rCRiUDopRWur3Zl/
mTktDRdrSMEcz2UW04DNxREpddVSFHpk7pyTGORTL0zg56E9alVFljM1/sfXU3NV
6vdOF3HOk+NLeDjHg7M5fGjs1+NojrrOxV5FUwuo77WTb5YYoI9c4uTykKzmxUEh
DoaHKpWE/HUQ4vFh+DH1/mKBu/B0wpzwSK6+sWtlzQPD64jqdh3phjWLifqtws+U
lo88kxuTfrcfmMA9jLbYN+dVoDNCKCr50sudpD9RdAGRoGAaElb0skX4jKlvUTF7
ykmWk011HXkPqBKDlnPxQN+ILmSTRH/OlbiuG5yk1mgsDl65ryZ6aCNZrXEKi6is
7JBcdpA+aRDfg8IvsfLmFHwJNDqrSnBbfcYexw68aKZS2ZTaZRuHMvxZy4EfqT70
tPlrVcXsSMYxS2cTXz6okCK8kKvOqDaPFwini2kxwTbjBrZyYFVqM/+8Fl+ffIRk
JumIuRDAbir6imSdHoWYGvY5Wd4fBKs15GjPBZS2qoWtnh9hasL4GJMKkhwV6tUm
aktz6/9k+asF/GxC69i4Fa4AMZ8yqmFzk7cy+QjSZAujJXpBxa4wWxBIN+g6L30/
1EH8GHqaPG5S1awz4nHwIHsSZitzFCYCZIGFJxUpGTlkl64OLVKFB1Fd5qu13oo3
qS/n0jENrbnHUnz6c0XzL963A+HZAbC0tQ/XiHskA3te+y9tSaoM+ZgFndgqLYIK
5XsNN9vr4SnNhv6gVpwoGdhKC938KfHqN4ceL3TrKs/kE0x+bwgHv/n5cSEDvdQV
uDUcc5C2O6nM840LgjE2N7k9hEUf33I0CqbkRWDzBlGKwRkuVnsdczwzakApRu/p
yDkiVlCjH1NPhKfhB0+DF0T0X8l9zilERa+/ayv7+n9ajPdTmULG/VoAh4ux9bUB
sJ59bjZaZCR8HzDXFVULsxDrZguV1uZpDwsybwQO2smfJJ+pKGtYddSx/UD1jyxo
JhhYJF3F6VqOahz/GkFxdYMo74KcxjwD3kbbBEP2N38H0wneNCgMffocRkUulQfM
d/yUWDelFmYm59Z2FCRqPMJYbxi6kN/PqilX5qkoGKVlNWkwHnkCxUz8MMJWnwJI
CPL5h3StYNYukxZfFxabOLk2jqBLiP9ssysRs294Fzf9m/s+AiXfQSiXoSi+lr/Q
ZoYTDN97Q1yhKOPrYJyXBt+S2KvUcM5TDil+f9MzA6geja/4qM5z3QAyIFnLgqFT
yUvVqDPalWl+UebSmRxzqGMTJsTEuJa1DmkVNiGfcs4B+817CshV/GYI1tizSuz9
Ws1vz3zFZOVFuhpvhinNpS5bOzsyq+phsX4wWDGzHFBfO+x7QbTs0sp2HQb7oFHn
bUWXwk9PrK+tU2lPeWERHD0ELY843U9uf5cowEhuUfbIFFx7sOTvn+jTiXxEWe5x
8v1YE6IvEmVdH+TcJ349FesdZuJany1dn1IajlDxdP2SM5taQ7uAI5VCNRGHzrY0
tvfKVD4jDcZ/uCgqIWwsnn4QgovHaT1GVEVUfNDIs2MjiSvjz9YKg7JXNplU0Euc
iGRYqXroh2GKp86eF2BA+RBbiKhKzM0fplPp4SM+ONGMDnQPU4W3snfnny5r30Ue
tb3t2zYPlnewwReo8Otxh4XO9KTeGTxrhEtw63kEfyqjO3fTa3wmET6igkHz0xcP
eIQtmc9ihuxfE2ujwM3WF0E8YoDrebS+EBFML4j4wETB2cSKHU36lbfBglc5FD0i
Yla6YfeNJPYXOkqSfpN6BVl/UNFBkqtAh2BRwKBo+n9BjEnhBaGJBThssmGD2o+4
mYdFMnD1iKq/tSHdrD/cBQWFEEa8mIlVlYIge4rHc3komfPdodnRsLll0gEUvDFK
gWoDGFCDH/5xY6ZSUztwKlKJxLXk2k1+UXtAcMIB/WNBwfjz+WevhuHy2dOXOSdQ
pXJhBKsvWHKGcbpuWHNuHPo5VP7bKhgaUZPdVzT6tE6d7XMYpB1b0w4vsyndBeE4
FaerBmLyGO2aiQJ7pDXmfjgxfA1fGOMaPQeIewasQI629OZftyboeMTIIC7uvKZR
L4pWZc4e5MBJ83dCBZfUIdX/WnQCJ795I30HesBPMcQok9tGDdgZ4xKaCNzwNifg
uAu8VvINR9pdbKuFv/xDnYOfCOhs9oT4oJ0tbzH2GJ4R5E9fOuJFjWVOYbWgVxb/
e3s8h5ayzgMPq8u6u0fE3e4I3k2VU6ZqnIZ/wmjLjzeojtcJqvKmN6HvtyUQjHP6
+96To4DYpTuNf+fDxMYiB+TKZqQJ5Z3ZtsqnIxlCaxvrPvvfBlBHfawSIW5nNkLl
ybg2vTYDGvyKE3D4FJveKqQ9kAOwBCtgcyr1t7ORtDs7jAgHMIQn3jVAq9oxcj+9
Hydj/BA/wrihRzc2OcWs7OzHL7+4UOuuBiUcrAoyuWLTHxphdLKEudL1AG3vzMy1
zkfGaowFe4iPsXWw3mfkZhUKQxbTGXwntpaELQV6puAQXP4irW/WN3XlF62hk9bn
SLzOjD4pvDkYKMtJh74GC2P7LOwpv9ZsRlU4U53Dm7GDBKVtVf7Vp+BHmxrATVPH
k37Hxkk5bukfn+lbWine0qhahUf30/JlIjcegHEe03zLsqpr96jfV1JSAxNdsUBW
zlGppA5EE45PdckuqVJxjiMmZxbjUAv4SScg4NiSCf4jeTak151PmQcYaT0SCV7K
EkR65rkA5bXlWRiCN9lrAoQSj9joJXm/E0ZuIFXG8tPVgn+0CMgdpnZZMJ8N469E
KwEyFsSMAFki1rDcxyZ1hDoxE5OkLtMKr4XUlaMpHa5tpnam1CFvfSwsqKqBqBk6
IESO4YtxqGO7CHmniVSKGn2R4mxn4QWpHU7pdJ0It8a5lJAzHrRSzKpBgknga0je
PosgYKBlPpm1YgMptX75TVqsbIvgUoebFHKm6xPwhQFhpakfd0D3Gxr6xLVgBI1i
0Kjc9q86wmY/SjEQwAuhHaoy/QoYyDmtao9kRmgd5g2fM7AsK+BR70cE5B/Amb9g
IVwqzNTAiDFI58zwQkQQL0IYEORxR6417Eg4moP3ZwWTsFGn7s32Jn7bwAz8ycSt
vLJRj8WL0vZuoGRU5o0exV9SP2bA2cH104e8rb6b6tSu12UJs9u4SD5c6c24lEJZ
IrqKg90wV7AEVwamhD3dHu7hAxyHkSImqVrFfo17+ltzengw+oT7KiRd/g4pdKTA
GdN81/+4jN/3EV2ppQr7lSLCOWg6WkNjZudUlZh+MZeQBd71MchZDNPDvg5DNifg
1zaLVuoVaor7Ydx7BHVGVc49ELatya3nvcLhdMVOlidomSs/RMQ5ykSMLsy7u0K4
BvspTzyf41TpPi2IFqIE1/0gLZi9gvwjOQba2q/5A46KpwBInCVPdtBIDun7p5qR
Ivst3ripTxdv/WczJUmu/PPAA2XJM1WMVJXL/6299blXbgKoqC5h5zzWjGBzB3gv
DiFZ0nxsLvZsWHUPp20ewzK07b38f/rZ5RG14Cam7gLPBqJRrLkl/pbLb9LV8R+W
omGIm4Ipj87Hm3/khU/8OEy/BUSc1ic3eJGarppu/u0FCYvySlbM5676xWdQvjSS
mTBgyHi799xR/niYzyDxk64c11QYZEYPHl+VS41G4SQ8oKa0cVw3y4cG3Wzl4ur3
wwUm+fXSNTHBDqBc2mxmUBBfsEpw2C83NiuDRxCYqI1cHVtDJ3b2tWqkDw68grJB
q37hqC+9MLW14OmKEJ1fSxwQvJz9AgD3KAbqAS2LmKSh1zcXUWgzNRkvDxwXNJfl
Ki38hLy3yaGHCwQWtM3whZIj11KBxXB13dKkb36s3sWYIIPAtaC8WDilBHnddg9V
/PzxLBdxxOFB4RC7gN2VCw0PFdiPBCCwVDabxXkusoz6V0SpQz8qG4+odyZwoieE
mfEvu/dka29jdnMevOXuvYPU/g1c0hVV67a7YCwXUMfLstpGYb+1k5bUiqQ1rQMv
BO6upDCXVjmahLLvYZcF+KC73LaM6HYazQLzBGeTcXhmFyzbv4NGfq4hx7ekD2EP
p1SC5tdnMrbId1cocJiT+bF1AlSLqOJRV01k9i+AqYwPzLUytfAWLqWkGljqEXEn
u4nEmbYbMSxgTadSrouIcRpTBX47sqAb+3N9oD7LuOlWqNMX0Eox3GbkQw2r24Ar
2GZs3hgs4ksm3gQUTRr1gv/sqMLk4gatZ0z1K1J0omnosrUCf8SI484iwb8DaqZe
XeE5AQDBs7WYIdj38B2fLmb7Ci0RRpRFgqPpazEav3C2H/AwZ8ClOIfWEHbvHFGI
YOztndxfLnn16XQkkLMx2wzU5CVUqqmirgf/ku9xU2q0F8QNdnE+TDlu0wFDtAZJ
zR3hH0gC3EaPbYwRvXVa13hgIvCqKGDgdPHy1rzH/RsV9P43ymhxldK+ijre+Q5a
KrOg05wsbAGfbnP0YzdXdtvJIuFoIYJkol/Mlurrz60j0bY1cPU6QL2jPI+kNDAr
8/jg0Lx8NLu8XCEC/Zq7Xt26QnkIjyisFsg1NnRmh+EvotKoQsKpJVnhM+vD9/Ce
bjUS8p6OWLPZToBRQJ0PQq5hAIKuWf/UvM1f2/+mCM4pp/9YuOmIVk6zsL9cJVrq
lhmNOk8NJemAUupm5xoMPAcm+t+q33kUBbIO+p6R1GzKoICXF3pcBDa5EYyrt66+
8crLbgE1j+E7uOCw1QSzKLpZJEXqLDTNDk/VjH8yr+dlQTYnEA+SeQWhU36bJE2F
HoLke+h4OXl0USa2B6IlHSaHxb4ailrjniliHqQTqG0K50j5b6twSuo1LW+8kVCU
Y5P2xk0nq/5otSUCNofADw1H2zdvPuiI8PP4MGgX99hBDXHhOvbUcb1FBzOKyPVT
SU9eye23KFDW63/Z2eRq4NAR9CuWj78X3Jm3izsctRTf1AjQ1oPGPflOQSgvTMqd
phmVNQmVqTI9w5mPanIr03rjjQOcAU1VtT+iQEwOlUJZBBjyFbfpg2pFpzXFawiT
2gXatu4YIMvwrbX/1iWiZWe8NYbcPORjrFC78pvXby1+NhNJiSyIdyEPN0wOWA8G
jGchQ6/rL3fAMQd51s3ZD02rIqlMAus5BNGNER0kloWRqt1kTBGvK4UuzpP3BdAo
28sl8Ws8SyO/PqnQvF+UCONTzPvqVu37MmrPjkcnQL9dX+Gl3ZLmugud9Dpdn0nS
/V31o7VpCiQ1TFD8GoLdBYgiYV35SO4i1beU89IZWSC49Tj+Y5bwfNWuzvkHKSv1
JNwTCJZnzYuu+pJr8lrjiSgNYdyZfWO3aK/wD3n92JDPClvj6e6S5u3KDyFv2Fvj
s6EfwqV71N0u+ax0Q9hyXfK7BI5csaay2s3judhJTycYYou65PLzZtXRX3wMa/70
tseSdGeZz/G3CADp8VlaSsFInBoAk5b1n/1jcwSn2k4bOlTHgP74Rk9q5IWMwM5k
b7PhmtHiKgiNfa8ixm4nZwCBK5j6uEIimouXEOnal0LnWmTEYWZTinn5qvcP+7jj
wJElGNh0w+oNdmyh5mk/A/DdmgVX2Bk+IFdoruoSUgaaQvXz1TeCDzjGntH2Hb3h
JHYrPURvS23BwvlOqSI28XV+OqnR11DM2cc+Ol0Ea2g3ebYj1I7e2t80zBrmvsri
h6/B5fJ86s3p2hMaex3mk5VG8xiMTsiHEQ3B6aFE2blcnrJv2Esz0mhpm8nP3cYX
q0KxM395zGFYdL3eylHhINryfBKX7Qso8g7IEE+L1U2fZY0RnI1ZLrp+XEVJzX/m
PBI0wutDu7NEACcbe15lI5VE/a2l/ERb7O+GGZBrYtPtZsqNJAWCHhGB6rUj2iiy
28xWBvUvx6p+Ay3Q9MdlKE4UDd7EX5Ev8ZO1xycttuslHhZdl9KZ4N/LQT3uVHYn
6v5+gipU1f7Uz9Ps5E+aGsZL+iznOgrn/ecCdhGkCwBUf04/MgtDsvwk6H0ocAtQ
kwxdpEnbraEg1Mv+e5ZxlhdharNHa8z06TBopIZ8dWGkz0fK80j1W6to7dXf9hpF
ZcAmOlzSqutYcxsn1WKs1apC/2qE4zCYAS8D3l7djJLGpzkjsnAyFaoTgBlq5mxH
Mi8VB+s0JU8tUjKgs1sXj7L9vgXa/AiFe89MDns4NtcZPD/K7QPETeO1wKs5gdWp
rogupRjZAeUsjpV+u3kMiKIFlo382+2O1WmKpwMg9sZI9HjyIMm0xD8hgHh+HLcw
zslGX6aizpFvghZ56vAlkYAGbHVrLV1pXGLvIkwY4hwKihlwc7w4W6rQpcMekw8N
2Fk5NnteFykcYcl8FbaS548VPg4NkEuqXbY11CbOyVNwS90FYkd3cgORHQihHmEx
C+8gBdekIMtWBc7XvXHxFvU92k/BAeIzzHSJCuOr1kl+c/XkYCiJapOYYOg1yqPR
pREY3Pw0xB3F7dcj2SRwFpv/qZcvX59y1iNJZhUPkOEQTHk8dHgwWQnUkpIUsvBD
uhYrKWbGoL1+Sm88MJWHoGagSDvG9/PBHFZ5/5ooiNhE/CnKKD6DHcgZESmIdPF9
uPNLHpeun6DAyuNnfbISBLQqgQ/gRshXr4ORA6D06C/tzbi/hIjo91uW8qJKdky9
7gqKqsWh9YaHZ9/RCOwSUra9wJc1dciNImNqqDjnKZ2KTOP0k0T5LFxSyZoUmUVo
7l+vR7mh/j3/6Ro9RpZl97EXQ2uVpHCpkVeLrgEd+HN02zNp8Y9KEnGjGnrGSHub
w/f4RLH3LOFOfcfFczO9CmmKkGgi74w3kdZNtRefDUDFzmc2a+7MyHQ26pVV5EgB
J1x4jeL57oj7FGFZSN7B2hcY0g2tde7SLL49X0eDDspEtonql9IQPYepuND2LghW
KS0BuLcshzGU6SQ4hOTdQTPgCx9KTlteB5BRUmP/2G10Q6oEs+n/FxWCArJ4hEsZ
Gpi56HOcejXOIvjZUI4LVP1f4HfSSrUY568z40D3erY1FP+GkBDUt3OIRE3svJJo
qBTDXaE5XIaDsVp5ScHGj39IJfP6flyJFXJt6wPhkGBHjZkFt6IDUFiblizQaXNY
vEI6UV7YGLvhpPQWsC2JyYWPJ76JtNXZuhT2DgQ742TDp9NKOZ7RfpGwdmaCKCbr
5WnkFiZmsgzXb+avr964IeKjaRyT+wTepVFBXcKbLdbvDCUSs2qQc9lyPwcOAAfw
h6VETIFtuAgYPWr8ky0RYjCQgj/Eqhiw+TuYdEwVAuoSYJbaQCiipFa3q6g6RpE5
dbDZfLAorq+3wif+QgPAy2Z5y15zzkJFNYzrLUwvYeeEhbE6QOP0vt6xQta5PiwR
grVjcXeTNeD6nHA9m3BKjfrJQK/p81YXZDVNVeAIYlAYYEtNGh3oBR90YRED333m
bvWdBh82hnPNtqaWmiuUvy5uV3JZbpgATIvHAR+/PXBxLoXM6XUFRnUcYED/lbz6
XHhc0e5Af/61bvDVrn8jYtUmO6//Y1AnXTWF+gFIwD1BjiqC0YnMmHMkjWJu75ES
L+4dbrsUmYVIv31GQgpKX6WPKBkXt/bcvbUctFfsc5kVBSBjDsGXl5lV2ygrXBUG
Dj/oPNyH3brx29s2e1XnHoX7J0ElADN5+zfhMR23+9aGpsGavY04lLMYi2KpPv6k
JAKo0oSWBmMsGwXP6KnrTf6JaRxvOvCfbuWQpGxFmL2GtdONFurI9r7ICKuginxP
SM51pvGZH0GSvqjl8xUzwvdsq+htzEfa9t1KduJMCC43YyxF59hK8rejr4zDPqlt
y7/72JT604ao+i7JF7tVYWQ9Mmeh1uCTASnn03EJ5W9FGdeuv3GUd1Y5txboYR1O
S2A5dpNUg9b6CTQoA4m+H6LQWkjdUimgOuViV9DGcQ8LbizZJhh8t8te6p4WQrCC
IxnhcBxQKTCNtwo2pYMLmxEVUso0iItQRDczbc7IFtMlZjdCTmS2aNtHV5BAQsTM
5sAan1iDpcAjXgjT1CfW2arj0n8M+r7Mc1fOMHz0pYyrBjibbCJUCuWTG+ssMqdP
iR8qT8hSuU71PmMdECg2K+lgRrMVwCJRqhocPj+sHEQdrkzM+9jmHekWbyLu4za/
yhVFuKtMowgjEZn2fAyrd/OgoOY5OV/u0Ofoz/kCh07ioGtRp9XwhdU5YQLijfcX
qoOqdZLlOpegqUb354wFFG8es9BUG0zANYHnvE3KD5qC/DqQnUbWSUMdEvbqM2jV
l+bh31sxRPuj7E0bQ02Au8KHQ9X/MKcSVGHNbxi+xloIjk/lgm4ZLsP0AybFxcY1
kfdg7PE5Mlc/IgaEjpDLnlhaMCwRTg9azeMJkEVpPS8ineL+mYqnJoG1elCpR4YH
xNCoi62xXZHsFhriTIgvgMcabC8iWhMRoXbAZ6JXIi0rVdqWUywz8t8njsuk/CDO
LKRvjztZQ4FsvRw2aBdZKaO1NbfPF34b2pb2ojmwcwbWRhOAmLd0pAkH1zv4mBPj
hsFv/98/Gm9CoQZtCOo6uJRjuD5zXt+65u+HaGymeCaWWPBUepdZ7vLl2tckzh2b
JoTm0kR9UIvXgMBqPX1N7esbgu/X1mqcQW6NQVkLZRu56YeTws8UDdIPEKESt2RT
hPox2Kgf6RAsK6BX8PyNZTbpuR9yQWnTqD+84dVM1gNdHV/BCCesLkwe+PKUgrh3
Oo3mbYQi9EzoOIfX2mXNovjmGil6iG8mDZArxYOLE21u/vN4cHrYuk/bpx8vDUpZ
L/7hFJ5azHK7xZjM+DSbyvWAlTnmLBJnZQCJB+SS91lk7tUFDPtc6azo57u7vjmc
lxXMNw1R2ya9TgCVubnmlu/pNfGZclvxCdkJBEAAjGMyJH40C4ZdyQMcmY0RIV2G
PyoVzjBTW7vKJPSa6/eiWl0F/lJXBu0WlZZk04F5bJfJcDlbKJ/zclft+DR51PaJ
XtX6Vz7fgp0NJ8rxrBP6ukPFb0V0WcfttpHose0MMacrRVl2lx7npFIRc/QOTAnS
28G2GHC0ANxnYtIjHebFhaQIeUaRSV2m8X9pCkD9uZl4QKVA8lioQiQgVEAkynUS
r/xNVq+iUaGwAfanz44iQqSCJg4MKJIfy9/HM6YzfuQZ7fXGYuKj0fAPhRH8hnUy
umzqh7Cc3JmXXN3e7gxsA97HAi6hssl2kk63rpeCmR9i0gy4LJSl4j+taApG0ol+
WGm7g3zs40fM9mJD9abc1664rqDKMago4TBaJEyJ3p2rs88SY8VujpgDU8uVlX/B
2qxoUR3n+cTJMRLH/SOlT17DfHRVm3E70LsQKDQ92Ah1oXZWN08Wp9Mx2W3aQ+cT
yHYyYRyFsVdK+E1QPZFgKOykm80wgvOYuVmsZfl59NZABb0RNyR/54uXObzqaS8V
y5Zdvj8s9qLVrXDGDF5/29EydkMk5g3f78wOMv1mfacyXeWuRF5xDtthaEoP5jQV
94dXmFwViAr30eXpmsKWrjK6IRtu2jiz4L1FGdO1dyP/FODw+trnwv7I+8yuo/S3
k3qCEVNHzWjxwO47I4iAcDYku8myOGw91888vOVboOboCagWwC8SE3J1izLAPZvM
gR+1kUTW+lKmZEwcdtjbb2AlltAF6TKHo/c9PXBEZmnM3btX6HovscpNW/eFAyI8
FL9OMMqXwqcHPWUEufAoavnovNHUhXnU3EqvcFpAT1MQHj6llhuTki9xiOOFPKyD
h3Tm1gQEn7ABfDh6G65tnWoTfoinGspRkb/tSeVY0E9ZKIq0FLb7V95o1TpoRxeh
yaqNNgdwzQG3iqL3V/9ZgxBQXNKLdH9Eb2SRp2uHuWNU3f+u91WQcnFVbIk6zZZW
zMciSMrNlBa8kXgqZIHTHfpFht+U9YQHklSg73brxpUrAuwuu/d0DlYQVEEpV6Y4
8J++62nQk8K/bHrfNY7eI4vdMRv+J6cQMB7aJqFGhdNqkkjqHmzYtqy1oUfOYQZ5
A18MOVfXr5aFJhmPl5YgFtdcEErn9RuV6nUsOnRkX8XncT/QZ6iBxQgTyXbP01Cr
kLzV+2M1IcZCzppvC2xjUKee8Un7eeZlMd5AUotNRkdoF8r3Yu72wZgejrkj2I82
VV4IM+xYvW9Xv3ialLblxdBmqOTZagkCGQbarUOZFdLr0lJCR1+jgQvzzD10uP2J
vvjeFhCK/tz9I3OSSH9f0Qu2TX2hDmKKJmjpgbbiHVcRFNdrIHCnP672fFvoTBcB
ga2FfArnDThu31L3n/iblfehgIYPll2IWso+gQjKdDi1tnOsV44vkVc75DdahwED
JHJe1H4KB/r8K91qWUGMUTjR6nJA/PpkzOW24TeEuVzT4VvXaGt1LH3Jy0bw9v3X
oSDyrecqVRRbe3W3Gvm/lwsUrPPYwM18NBMbHF05PfumExS5lKjRRvY0E5/kTglU
z2Pqa3D76Jjj9KtIZTB6F5TbqRllMsDCVX/wkr6f4RtdZxe67xDSu/4QVTPEOqDx
KE2LM8UwWY6XD5krqiDXWik74ZCN8wztgHXBdniM+fbYS4GL4mX3ShZZb2oTO2EJ
qKrxJDjZbmh+y5oaU2eyqedbIgGDZcdBs4Ktlupj/Aj//zKDi3OntHJB/3gyf97U
iWlYe21MAW0UMkcwQxSFe4QpidD5sEDwTSWbdc6n6CXU8aTRgxRGipzD7ZnJ03Mo
RjTgnHf24Ig9nGix25hF9VDn9r2zFLc9yDrHWW8wYFQXK0ptCybMsDu/aIoS4M0F
eQxF6UkrR3X9JADWOubXJHfyh5H0korNtKTUDb9nja2BaniDGvblDFu+67457R7k
TwDih0UsJ/YWhSHPEiJPcE+D7sK6KOtK7EQkMSlmGBmzoZxeJFscxvGWVa+5pJTs
3rnM9AYrSfeDNTe5cIciJ1RS554xc6QBScgfPvCsMHvmVQ3Op+kbvjmLBbCeLwH2
YFoty1kdERyb4knvRmhLyNOtXy7FkKSDAc6jbK46DuYbSXCsc0Ros/3+BsWchm9J
khY/1q9m4+LiPAvofkp56kyKU8Qed4N0ndBFW7cy6uVwGHXNSpCU9gNZa619rZ+d
UQITsG4kUy+LQ6623lJaKhHDv4edo8Jom9dp0AIuKB/FlhJqLMXn6i0wVjtDOGCM
89RTw5PytU1eVSXtmPGLIgKmn2WLjNaQvVA2pM6XN1+JlLOksLHbsmajQkC8c0oc
LMKBsny1CfLCNEdr8ZJyNkAgVAp0UocaMy5VJ+WHIxvQBKIg4mrOld9nZYcoW1jl
SeeEFmQ73S1W9M1U5MO1NXd44UwmctFqVNNHq6bo3wXSSy7NWXaKgBbvhemFWPEy
cL+4I1u/MesPmfbRPSBxH7rR3dhdfo8Oz7QMgqS9MK3e6BZwdynkgTe/V3ZFYhCm
/pb+uaL8Q62LAZlf+D9tI2qjNqBRs98k4jwNWHXVyBJXgYo7v/0D7AF42DJjXOKD
zvz0tAbTJRbXoR5S2FNKEaFRb3T5Be5KgfrgYvqE2bGA5Rsv3j3WVoUkhKoonYRT
GZPeYZQM542tER+nbcTPtRFXFo407dIBBLviMzsV+z66I2Jisya4vzU1MYth4D4L
obAT7LFnwoL0jvA7ZrpR1zNH47azxAvHwzpl1pqLQpFfP8xtBGJ9y0nCtS/Q0Iyw
J809qargOJluYD5rm1XRblOZBBYFveyYFt1m0aIRYEexKQz1AGLVclG1NTbugP3i
CFGtNvNRatZsXWVg+pH3cT0wl+Y5IHFHId6+yt3Mc7VCgY5K3L0vHv6fwrlj45rS
A7ohS2duG2w/hoM7KK+pu0/F9dSlq8ScM9jKS+/6+IpRXx2+prHuEQxXox9JNdb+
xMulCQvuvV5Ix6vFMFGzsyR/jjPyxq59Y/B1qdsyQN6WMtA+3vlHKfxaHNqTqVTi
DNJRT/JN9bHJJ0ll4IfGJz04Kcw+vkWLYfF4ZA2uFgNIWxyAAOeyci5KBS65THyj
MjTMegTpJnEkIfvyWtTo/dzIB1zj7j+2mYcX3qYCqjr7G2bj8MbWq/v7qW+yZfkH
Khu1QxJ+wnxbpMNIpewauZkK2Ju6TJsbm5y0OPh47+cH55Dyll67B3dRXy1LZxxN
AYFQpXP1fK/psgODKOwFSdZie/4qleSOxrJnreUZ7rE/S7OlyJMoNrEaD1hjOluO
CYr+JM0xBYv7r4YQrt1LSi444oexv4ScVBIp8aI5hP20c6D/UYwqpPVgZE0/oCcx
CpDFf9ne5iaocoj3Sjbj86ou0TCegh74psoPibFCCZplhHdUY5YOWef0d77IEHFj
avvoRmc9c8Qn4xpe+4HQVuVd4URYw2iF0BXFo9E03IrykzJJMS72sj9I/iT7g6e/
aviV0CqjR5bPVt6+geITSvtcz27MAFilHfssEifRRLWnCyNXNN9Ykhp9deMXIeG1
H+1wyXxeOyPpVhq8FddS1JyZJ0b/U+YkDPwq/bCIRUAcb+gYOTqkSzdtpDXFoVyG
QsauIkx5Nyz484NBvrS1/a8CSX81Qk2EwVqINRUHHAq1Ewd/VVTy2wzvvrl3vFr7
oTcfQVyMEMHSUWtMLdOEeHfMR/Pac51IKySRhzkcQwQFPj6LiJ/vGZM+SUcg4wgY
xsgFrr3yjm5rFBsIfaEca44R0ImoA0X5oOe3s5v7KwVgtJAZiGFkBaU/zMaX2irP
o8fFE3kj/xWaPAOpEqEA+MZQvYZ9CPgnAvejXyRZuvOP2FUq+gIfMKnHhHhvF8yv
D1ZJm1BTMT0mkljN+zJ3n0xUyU9bS9glxS5g72hfDOhDBtSqeMitYzBRvvtS4Q4E
doyi/3+F1La3Uv7k35DL6cAHhjdaKt/HWTnMRmX1lxkSOJrcXaFgttgmqvm4gEAS
2qvR/ph6ablhGiQcevsD1mn/PI9Hr+0zaBKJPUeDeZ37ewSlCx+bQSvO7R+2vsCZ
3AkRrZBV4StLJ/MeTNIfc3nbpbJtVxLAWI7GJKyZP4RzQbnvxEIZ3V8If/eWJd0W
pd/E8t0pmjrC6JWxN3h9P5iImcm28iHBFTOVJoBeyJobN2ErS/oxu+6j+3SE8l36
YZoD8lzvC4FEtB6BYEeTs3/Ht+A5aLsl5Jwbhoe68a7/CCmaMSlbkmBB+qIW/s1e
6erPKNFRwONOT7Jd0FjyGpEGfDtl3v8SofEn9HOUiXDbBLFx5YbWGGIn0fCDw5iG
dP07KtQG70d4bm+JXjWRoqKBj5+Ia3g7DI/5SrxYLFJ61a6xy2g8aIeQ566uHfFF
B/mWGSID/AzJz3SzXXsD0Dely37Rf69ewjWmBuyBUqJGslh4AC009BveEnRdKEWr
MoGPwHPxyT26HYX6pnjmpFZuAPDgJpc/XxpQ1zHSnih/sQoLPQpngwyWsPqFpfNn
ZdbBClhmpP+aQIWMA5gSvQLT489HaquBFrLXBdoOAY0aIhbxgeJLoHW/AraYFlUX
z9LMoTD1lUjCsljbSfDUKSQbx7EJdyE6a9hNih8v7Kf1iQRE/ePLlABZbFAMpRdy
bseWrXiKxlMw1si3Af5USSE0LrXe6czk14824qe8lvZx7y5MvwZZX6vh/QkkWrGW
RX8QgCL6WANsiEmKQLZqRC5b5BW0kUVDOutJJCnU+xPcss8sQl7PzQHeaPY5gL/Q
eze8TwX9zWemxri5gjywTNk5qR1fY0MGEx/TiFcTbwmg5IhTqCR0bOHakBG4wL/5
AgI0/lu1tvhoDW/Qsh66WFxqtNpRk9GTbzvSub/MDlwhlVwwzistsqkioyjMfkX8
pqBXbv6kNBgW3KBZXjLI6nnBcx8U9m+4EK1L5ZroJjNVQoPUSx1GmWadNZ1EHAGW
nf8wmsOfNxu3du57E7yBkVvL4SsJDORal0CUs7/QMXGDsS712/gJ4lSh1OPPgA5J
dTxju0pNd4xffELibXFXQCaMKnTTJHBhI8Es7EKvIChYwz3a1f1UiAKOPMtqq/O3
a3p6r7Gkee3quW3f8KbKwvZwaQyjHWcGLxpJjfxhegiPLVmwbFUQf6M2CCHYgvEs
SDDhr/VPJ8JbRGic0Dc6OMi4sEfh9gsVFogvjIBxKiV9RCaONU2HeZd3b+bvy+9n
YYTtpaf9R6pyhhQWmlUI0Y1DQuf/jyxUFJMG9eWxD/EUjruBE2bErNVaJFSyu1Dv
d/8vMmM6I8pXeLzzJCJO5Ano5OuV+P1pH9DsKGMG+jPYJlhlKOsrvttg1nSyzbPR
GwZDTlURqqVpcXgelhJS8OOiFl3JuBo419Idb6+fZksmBwxPo05bBdfXYHeYAYeM
mEKfh49cLES4weUUyVO/BF1EIg8ihesulfBdXiUga/OA+IyR8BZ4xFuOwGB0Rajw
9n6xuCQkcRHqvHAJ562Or4NX417UjJYbmcoZmHk+m/qDNNFdu81D6oohfvR2+Ehl
wYw+shLSCZxveudbVq1VR2K4p2tFTLA94ltLd4YGbGq0BJXZi4/QTGFnlwVEn28x
3uFi+TjD6kaAKuNPcgcKenn+q35wjps35Rp3ShmJUuttEs2cw0ZVcd1biQuHRXNa
WVL1sT0L/XTQTCecSseDfNiIh1dwn0mC5WbZX50nz7lE0QxpDsYXDa7D6K0zs/Qv
c0Ik63hPZl33jXnquFUqt01/Yigl8aR4wabBhFbJV3kCVp5LwJmUgMR7U39d3kW2
ZUVGEtTBU1cQVVbRHomoTpaN7inw9HZP0uQFmGkTKbrdbbmTiP2MsJbHTbpDqquU
pDE+M3I2QGyfEqeWTMcINtO2Bdq3rHs0NVt2eWsrlSOEzpNGKDuWCUs+K8PtOjGW
uykiLf0CVjXz7eAdFcgQPQ8ShMcAU/981jfHscJWVLflov3oDmRsXewotyD/Wb3z
V3UOIqqCB3mzfTFIfeXO/7W4SUfmdxh+CGM58Alaq87ApR+fEAxRX9jNUWPOT2tJ
EUGcDI4hdBAFES2dTwUT5gP4ZPf3W42L3bfMbTm76qcn6n4CcaeWj4cUeOBKtewk
MB7eLkEbRHbZpMeU7YwskcDgtJWR+dLpm3tSEOjlFpiQPDkKN8OsH2qRgKo0+F5J
xK1BozvoAHG9AsoBvEPDzJu/5N/zRwJdtkYkGCZFRq22I2odRxQVLGc8TxFLQqhq
aLLCQrwKOna0walttfXY1cJyMnh/qZBMF42iptIZp5aJAYWWI/ip/ZCh+x+0Wjz+
2bgur4A4TksR+UXYwUCirWjlMu1WPak9EieV5wM3aPe4JiUNSehYZuVOPdwcMO1x
th0lRpn0H2MEjQ4EbUMJ0Hm5VaKTz8bv+YZV1Kfx5g3NUPxXFYdN7Y4ACWgNWU9G
KoAPznqxRMtx40RBv0Xg3SehRCHdZM4Lz9LEwOwtELk1P4ztznxTfCRqm8ASzvq3
2pr2RDxVZ3nceSlv62RE0B7Xe5+y+IccigEuyFGO/mYlQTBXI39wj776hxt6zcHc
zmRPF6Y0ukKKBmEiIdwaTj6bZWKxWq0V0mEfBJW4vE9qxK7BL/UR+eXgckwrLmQQ
t7XrZpKkDjTs56Hv5PKsHmSZiZaJZvWHGeQUhOSTH+BHWTZcalhnuRukyMAh1NcB
xdFihZ5g1rKn/TIoYELZ8NwGmSCH1uKgM/f+o+okTbe5Ckww6WYroFRf76rcC5UF
6a9ALK0TfhsFFcu7qPzS3c4/mk+cjT2A+pIaiZDeZ/Uje9zQ8ZoRsD+C4CSqTmDa
8/mUFfTYkj3yD+M5cuVxugSd3zmWfe3Q1+kfmj9wpC5/fH4nRf5Tq6mUqEGN4iC9
riUpbIua3JzonQJz8MZidM5ZwUzY1aU+rGL+olwJypTsaRoQ2zAEWf0fz85D9qcI
cXR5GZ0TAYoO5pkORTJhLSTaL0RcfRSQYaVV1qR59zBPKX4lD8CvLKEEoOcH3+wK
8sGI/6IEW0kfKzaNFJYipLvBhdsBqPMsZJeFDlyrW+oiwXsW4y1FVGZCw1StUq/C
eZw2nfZK8NUHMGwdDqh88FBp6XQiR7aETT3I3tJvJIS8SueyICSVaua3n5aUKTnX
sPsesYHQMpOC8jbrVAzocdxKS3ZBx1gsZAef0ysnxkWKfzb9N+psGgSDpdp1cWt3
bhL5jU82V+zqUf/F+O0zw82TF87D/k9i9GqTuFucp//scXnSjPFeMu5husaCHOD0
fqIK59dgtSC3y8SzsawulkI1Run05OE41nni0PSK0cioqDZiHvf53vZCJRBhHJlC
6j6OeRzcAo4Y43M00E82nImbuMvRfl402TvUgncsWjxQmEFUxNOySEz9+KCtHkTb
azD3s6It20j9P/YsJox8+/4sRE//kKszfs+q+u4rxRzsEXSoikAWNGLq9PIcQDs3
T8LpMZ9FauI0RXVGPTDoycJj2d5W4AJkNn9aZ5nZmOHzXV+dDacGtQX9shUC6FhY
TV9dBad1xG/r0agZFv1zt6/em3gpgJ0mEvd9jH+lVYjqp6xUaV1Mwa0M+4iJ+CpO
rOfbVojf9l3tvP88S2h4FMrh8YYSPxPh3gLObKcZznRmmfkClxsdG9KAwrhwafsY
UqP8u30wkEjihALjsOW5oDC5YI5cMd4h039GIEeYp6D9bU624YLWzWTTEBFYhRPF
TV56u41pGwkqqBDTe6seGyf+pKEQeYvx9jPSTU+px8uM6jMvBvbaa/BRiGD/B8RY
goxV+FMBBuW+GwMiqypPaRhswQANVsOn02VkvvmZFOd5ZKG15b419vSxM3xaBpyJ
OQHj0aK6uTUWQk8BTPiQ8U3mg5W88hoOpolNaXlzd1iMiVAQDttvJR7UeM9LYWYk
f9tjvhtOW+CV5dyFAVsG0YM8QsgbPDiVzi7CgTeBa3ABdnG4Pi7XkBP76gYWpoAQ
VxK9OgD7bT5aVFaVNtF0xF0e2z/9T+69hAGUc3ZVnPBNqEcSyfdp4N3bIf9PY0/l
zQCTIXPR9tWvoTT9RehedQgImI6jfOPSUtkwvQ656AejhvZQ/Mzk4Y/SPWNF1zsb
SvzHSmG3U4ZMWjqCYWEGozs5Grl0KuxgEhiegjyq4XYMD/KBgDgAnWD0C49BjqTO
SZpv7wzg/QRWhBBZ0Q7KWXbjtQRXGxZyOuLUV11CVlZXHRm7DXeeGqDuqW7Rq69a
FwJdfrevvIJan/zY2TklQUeGJCIDmG1zi4ktfA4Rj9scFety0EjQv0rONVBd0zIw
QPv7AQ8YYFJX0S29ItD1cBGStlIZsMYwA0u6bGV4IvK//R1EIeey1814dCtyqO75
AUOAPqErc8aYpJfdC/Qhr9wAxWGlKZ709en/fGQ/bJWtYFvsvebgDyzg+noWbkkO
3bMUIhPeRAF/wbUJUaFXuPlFFDvhNiTNAzgf41KR2S8ZkE3065Elv+A7/lWpkykT
9z9VudvWj+Ka8oPKsAcayH4ZBl7nkhEcQ+7ky8lFS/3JJaspGbfm7dG3UItyr1pF
lLlb+65m3hV4DQssLb6YU6ipymCipstnWSiO4Xefi6xrufTEzeZUUwrQ/T7s4WGj
nz3jkVlZrBZsfSENUqPdOyJGIWsq6NCaiSX0hjJurim8RKlGo4p4g807g41Z+SpP
ErRri3zIzPiG2bEDHa5AZxlWEX2GFrtXf43vBuPeTuXCA5nCd0oI0s1qKyZLaOJb
nW2PE13JE2t2//dDbpgEXqGRfrrK8NyPuBY/R0SuSaUTYsuTNR69ZTBul3dLHkS/
hkVjUOMrrKwCo3eln8tJSJZfywZjDvyPa6Zi7E/Six6uMFZKpROtn0E73Cn+mZFe
uP2//VbtJKyrsUi32V+3XWQlRFG4ylrGcmHz5sGyAGE/jAGFFTOiNlql5qgFd7Mp
o32a1VbjB/gOOsBoSrugvuEn+e8x//oy7XGTLzKsxQJh9a+YmYSikJlxwPm3kBNa
sIVbOQo0Z6GVneyY9fEDqP4q1I+kedZcnwQ/HsPUch34vCCvRSIRQ32QxWyx1TiR
8C5ycs+qXi4RVy/0b7KKnpgQqOJo5gK2YQMXFpxBVYFauBug32yU7dvPwa1XcPEf
5HLrNC8fkmD1gp1in8cxxJ/Qz8LJSCaa0yjTE6fCl3eNcey+5dRUkuAFrFu3VUnK
7FY6fiPrrHLmIjS6zSKcnkMn2kgTdbiBQT/RMbCgxAofFh33JfbWXWOPf3CrS+z5
8gEoY3u9q2Td7o0hYGTKiXQFnsFOiiD/wGZonIHSd4G68KYFY/5gTUa7cGBBQDMo
adD+Cu8w0ygYDiyBXs7JFlKAs8T+PtbDBlu2/GSmWiFm/ib7IN3+7WTroAgNbrMY
obZyZI4qAfjsAywQnuj5L3ldwCUmHAR2rwdUIcw9wwGWxbjB2+f/GFpgND9eDFMn
B9Fyq/VX2CU0KPvwhirnDoz5CPG4R/98hKDw52ql1If35/mMO5EC3+vcJgBD3XPu
8cs0w2vsEyN22GjG539Mqz6YCh8868jtGm291lzQXU60oJdxyd8lY/MGo8aQCF2f
YYEMwFlujqLgWSFogxdySTDqJjFDtGX1WZIGZEyjGLDWepS3UQuZcHRkc8F2w5sX
01ZB8rQJLJjPRlBwpMR4jd6QyltTMAQ2v5YHTuHzNOHXnOh3diNXAitg4E1yC7i+
AWkZgITeQH9VKLr1NsqEU2Y9zpivdEQlUzVDmNtHoT22CxI+nplzBjgF5TyHvDhD
UnQrgYR11s5P1cx3DI951jHlJHpB0+JbAAQ7TAenhiAyrg5ueJyTjkSLFONbYQYt
8SKbmsofTk0P3BPvh48xjpYSJEC/v/COk+JP+x47ISHLPd6IvoYxx0fz4DKWUDzk
wNFbtuPLEDN1ncKz0VinuKn/wtRj8+DczMEQLJ5tituzlLlJiumKJ0Bx4XeaFETs
RrWQXXnd/8Kkuh8FotyBLkCUozg6yd2xqPvXl/ErNfpWF74cdPgBOo3j8XNLUyxk
6lw67znSmuJhVsFV+O0ukJgUZEcLaZgzmlayN0yVkiU2EfOeCeVU9Ty90pYv9+Oj
5B6hYUtwBU9ZbwBDVL8aSai/KsDQY/aE9saqdl95NMqlKt0ajhG8x1Do2kxNLqCz
JyejNFHfsA6yUZGWwSJgiArT6e8dJOJIagxJxAICG3VpmxAVbUNTaBU+stcIikwg
4PydBPxM62OMcLJ7aGgK3CFNpSaSUXRdehzs3cmhy2nagk8p3LfEZEfnhOBGt5so
Fi3T5owNQB8/Yv0hyFmQHfCboSHSbmm2RFpyIYWpgx/pDofYFlq20kKj11leJy05
VVwVlU3EYL6zqjAnzGh+t9EX6+RVeNpMxdLP6u4fMS4iKrAxMY/1jj3P1zYNZoZK
AN0xGvAspB912GXCTMJDyGSpqMVAYR0Bv6jLqfP658p65lnKLLmSCpnh/xOZpfRm
x6fk5gOGAWSkDHndWLG/95c5IxzwWGJKkzZLLW4oA/Q/upLaKdN6rsT9Em1YtezY
/cTJ592M/VWfxgwuypph8YpazSRPHnmUSemlZywIZE7zFeX2frDzFrA4cg3DZcHN
MrPkcr6rI5zXH3izb7Cdq2uT30408Y001wU2jaTRgFgRPU9JWJg+gzSIQTFLfxDO
MqdunWcPkGVj1IC6+M5unrS32z9Ec0ffmnEG4E5n7IAE5Fl/yGn41a3TPPDX6U1v
HCQFcSNPY0jkzwEFiwSh7+Ip54GRfOO2+yT3fACYi02jEX+U3AqFWdA+GPUv7lqk
X4xQHIcXGzEUMOhdD7fG4y+lcmni3PhLAzjLS+uUZ6A8J8YaFVmzktgaR79DQN6U
DSWRI89n6+cePWwWtfu8C1jv9IpyF8OrYqqFs4pA8LgKxPl8U0fXTHLX75Jn8PS7
dz10Jl3wQOn4oCxUTgm2IS1/tYIu1kByNNop+hXccZwtVGppZDaCw2sLC6ZkWTpC
cg6ndDxt8nGHXhHgUFgYbamSUhF85k8hP8ZiZyYNRNXMs95/7c0/GFH1gLK9g8ZX
eKINOJuyutbrvM5qYd4RUQOFGdYplEqYD0WJEeu5HWObDAxmTh0KAfwHzNy4Yj2+
UwEPyigj5tY04r1VV0SdDCy+NETJye29A+f5ao1b/eVDZoCv1aKw1E1BFdApP+Io
VvNiw8PEXxdWRq+M79jF74Tib1UhP6n3/FpsgWz5uID1BtqZ0ztwtoeqKwHuNaTX
dS2DhoykgJP18NxX1mS+XDimEDLAc8A9tgpml5zablSvTpYsycPXOYk/p0toK5eV
F1+Rgm2lwoysCJQirMCGeXGPc/A6GBGjPcHxMIWEl4vK2YOQuHrLNG3XlhP4G7C8
l1cdoX+Y0LEHBlTLdxSM5YfVRtFc1C/xAp340U1UCA11NXE7OXDudp8ZVFS7EQSv
D8hnbFUpqC3JEIc8iYKG4HJgve4hQEcHu6U0mba2fzrrBKba8IsNShGCm6iR5MhC
V6EorQ9wIZNP2krbNSG1I1voQf73CdSbqS2SBF7oyt8DTcWc91xHXeuxWgksuJ3/
uG7SZnYYmECeD0rLRUmO06kkY/NCiIOzZpStT7/jgy26zPP6umvCTXiI0Ae5Xmjl
5b0kQ2XRA23mMVnDaOSc8XuBZgraaU5/yGBSbd6YbRNwhjQpqPB5II2jocVdAjr5
qMU+C0RtlNHSs1XdT6IABGXGqzvupmS2EHwvEQZEWfw2x2fUXW2oveRewlPzB2IL
omTLLKC0IkVdcc+VdeJZc01k+juOHqWIyckpGQHEv982UQxx3+vcO2ABsyF+4K6/
ExYVyYHiEemazMqSvoT8QzjYwwg+kCX/rHhK23FR3cptZYVGEHprKuIZbCsFr8en
bmAzZ1B3lp5Tdhx99IrR43izYCvOvnYJQuYQpx/BmPBY1exZmXvYcsiTIpOQD9Mb
+RplOytJpqPJiRz1qVBqm2GcBdelX7C8ZivurWw8rukaG2MRBCscem4qs8p4DKNB
CwIQCkpIpuw/TQjkOYesyyUO8Smhj0wZ7IZe+6eWBJ/VraXCFqSNv1ItT0g2y5gJ
YABKaUGwBEd9+9knGYSqox3EAaPsd705xZsHwxvAwfapcIioumqFgu7dQZHiDFy9
TfAtbN0sV3dDEQ5UYsduk9BxXc50b7yO8+/GRPnP9VDGw1m5OgQzp+xLzAnz5gS+
gBsSA1w31RBSWHzI+HKP6SQsH8ULv3osgMNtEqAyx536hRtTqtpw4ZokglXdSmrq
uCZLU4SZi14ZFFsPu040krKcypyAnwPbEw2UkMtenU2AiAQrEfyur3fYL9hY5WP4
egi5n9vzlUpLv6FJ+5iZpAI/Sy47h+k9smhEhPs/6lb1F1vZwfwaOF+DRKOxlyv3
1OrXlBbz4An4L2TcTWemx/rKsinMhAfC2KpcaBDibwb+8fxog/mtZf6pvvML9rjz
qBmjp8Mi/y66j5Fw/GiBF81/9mQ57lonKds0oVTLRHbyuKmnsI1yERktoPgvQtnH
1qP7RdVNMYMKoLRtLxmeBLuUAUe3+C5ZX/XJRUqebQPRrbJNH+z/0Iu5za6D+5+7
sMnHdUsGtLtgpCXmCuLwz0XQUblEQEMqlde/Uh+RcxbhY8PznsyInNb9K/c88S4+
20PDA7d1ODw6Hn2glzCCohuoDt/gT6nC1cOf7CI9uUeDy1Bc0hJ5Nf8VHCCHfFum
z8MmbAtBy0WCmsW/QRtyUzeNz1uzL/Q52IvMcckyEe77Rt3mfutLyAMkUYMHvfF+
XNwmlK5Gj6nP1HyD+7lwS/jX1LbqNL86L2BqpoBsrnfxlMoYz62vyGVvhRmBdLKg
Qzf/4yUEmMJm3RJn8c63xcsZPgB9zk/mVdr9NCEabReVRHUf6vht6383UJVT7N1B
1bS5oSMZTgGa7AOA8LCEQncEuUdPlFrAS6nnOmK4VX2I0Dm4kYIHjwwc9qXWQyDZ
tdZid+CvEj0pVSGOL0ZLr5hOIsMoU5Jv1D9O0CNI9Dw5+moK/KlFydZbtUjOlX6j
3aZ4evmb9YrponfiVwe/RaBhqAJmTfaePIBqUEa3PjiuRbn/oL/Jo0d/SbUqtaqU
IAic06zgIhRZfu7H/YjazbJU+LUDcM2Z9hbZ5433Bd315svlKCAAtCMnNmi2Kw5r
xJbh3kHhT/IGTHn4FEoU5mR96Gpi9o8gYhx3gZrmEMhYyn0b8Dqp4jJjGk33Dd7k
NO3d+8uFkW//Z1au+Nli28mQYDuom05rbsXTgiDsHH/Qibepc7lmmbL2BaJKNr7w
WM5WziteGWVHlaFB0why9dPczv9bm+cioV9g4Br12gefNqAAqNbSOnFEqdjgbhIg
81lC/QZWG3xtvFMD4woNqYyxWeJls7VmOOBD4dhq8leqZ4qosf8yAPToQEFSOfC9
m1lT1F2BvRFkd6WhaD9BdBlounFwGUK2FU283HuCD0yDUXU8tDJ/MUQ7ROvMwxWH
rYexbSYxfgpPO8HwvYkzl2mPIl3RUNjHgdwUlCs/jyRRuKqu/3cwEiLpdoy/XMva
t1h1GtfWKodJJsSL9SF3gWTp0lhi7Ufvd3N5FfwHS7+eQEBWYzJ91hQPHRYQXclL
0iFDw2d++spk1MWccjyRVK178b95duAZDq24KR1qLYzh2ArPvMgj4BG5F2H6AjU5
xit4hzv95zmAQpTFl+gxgvixyZIMydFhWrW4+we31QgInWrb2oZZJbpk3pCOj7Tu
7bRMgMl28XWSvihyiV1rlEwnJINBDMit24mOVCPKmuws6d4uZAB7m1I3BaJOy2ku
aZwa6JUKoKlPYc9ttL5U3QTqFqdixcJbhu5Wy1e/Eu+ZHyVpCvSbRZRrVyDR3AbT
qi69CdPxa+lYf1f4yMLkw4dvHh60OJZvZU3v6pvmeqGMTm4IGiDA0u7ZHrMFi6Lq
04CfdE0mJ6j9rKwok1nkK7zbsmN20u0K+6DskH01B8w17qeXSTjtbQax2p33zBhr
GDTct1x6gg/uDwPTnJebUzRu4bnkQGnUDGgXDInesJ8lwbcXw6ydhW8OuJkEh5jK
sUwvy0Enmml79F3emQIwTDI6KU36mKNK/HECOtYHyPCPuUX+5Ue5VvGpJmyce14Q
D0qQGJ9cAm5a2bT1kqNfoIyYdT9W6HwBhHWFU2415hiD9hARFWYJVPxj/IjKRMdh
wUiiNEziAZk9MBzTSJBQMirT8MV4uar/pivDWdyWVYY7xX5NAzXnEyt79mtIfn9c
3LiJQSUDeDYXDHHOgp/ft5HPrIEppN5EF6PKoH62GfEibollJLwuTCbponwvjyre
7RxdEJwo7+YcEBDyoPckjmGZDgsXJWI2Bnk7/E0foSOCRK1aiFyeXdDOpp/hmyCp
BL0Xc4czT9YyjGLc0Lj+7lfAKIgZaw77zFfkVUtGw8l+sMP03P6IXyawbiKXlZ+G
xhS9JN+VPPFTFThE06PIzIaB7TDF17bbKWDPjMkR6spWevkks4k4XqzwL6DHNNZq
Oyy04kA6ZI8kRIIhrglvH4CZaBZvBoDng5oWuG1/2OGsAxrIeMBBNxmoIlLZ0wjj
Sb0rGj11WHtdpipMUAqXeq5IBkZPGTBFdgSMnXVknDDBNsivK/DnMXmAYTxER/ZN
u04Hj74L940Ty/kfdSjK6g/Z1XKWbQvXw3ijQEU0beV3UonaMqz/gi2hWErzTlf+
JveDUo7a1AVwIeW5KoZT0BZRP3B/P9XXEyti+XV5Kz09/q05FsrXuxkgZn5Kiip/
ZKdavqo2zcz+mU0yu72IUVdrFom5HjloHepBH/evHU/FOtTaQA1aeIzH7VPQ5NXw
1xf1Qq0ZEWLWeaM0n97oquH53fA25IqZ5gGYQaaZ7pHUo99UwmWZR2Jkg+/cJLTs
jl8tAY1VTBuxKgwjWfQW4AY4IrBgA+xTA8Bi3LC0QJQYcr07EWn+iURLf7ovEUwg
iLZCMzTQCIRjbGHmQmvcO8BLaGPuUtPygFOk4zRsjfufQoQYFoMap+T13JJoAE/M
z/Pqld6kG6v69BHQF8b5Dxbap3DNPwXArIw/sCSrTgIEYawzmlaps6W3azZEZrBC
OTxG12Iy1jO3dDGaXbFTy40VFofKABjc3pcI5l6VBMZ7S2j5eaXOVQq+G5udrJTm
kOCIt8kfAdV3jvOsSg/ikdmpOr4N5ZqWdyAQdZ8d3dYtxxh2vHNkrM19Rad/+2n6
BFyApkw70PPivDuylfPxDSzWR23zGXd6ICXa1nWrst6PzokZVh5PR7RYhmgGlQwF
+0L3+Y4N/GP1brc3PnxpB/uoN+0gVYUdEJYOQvEMAvbhJpChSg771ofM7TOxcjCS
TCNWZKp9ZqvUTF8T7vcXfbo4taWxziJZC1GT+h5b52kZrCwuO1pGTdYmtiFvqoWu
hePJDR+NNeVWDGkTBmCWkDXaueuC8QZ+mZUhB208DGxMYDCZGkLvjhBYvnXytyQj
E3CtQAv1qbya79V2T1Y21aGWyGQY+iK6JlKt91TOGcmHZUgcSumfM3mXxIbFQYh8
t2O59yhTIk7yeC9bMnq93ymTyZnrye37goldHGPlsAs03vvE24I5wC7lU98xqbuQ
o5IyahQA+Ce3tqN/3OsuV6NqhEOhL04zu45pRAyg5mFQADVyP/lXik2EPOY7O/5G
EJpm2+ut1+ybNNG+Zrvft7+GUzqXJ6IU8YcnV7eIB3dZs1ApDxCJoh3g49LEG3LV
ahoJ/ABjrC8GZCW6fwH7gHaOMKGzpWi0lePx+rQhqVDxGrlv/EUWvzFflotzRQDJ
Io5wDrebdwnb7kbxWQAJRZTfOAPQ50cVzvBFZwEesY9Vi8by0Eh5ufTkJXObjYbA
aTdEg5mshf0YQg/wJk/dvbZ1g1BZ0RnBXxbrcwU/qhZ6LbE88pCGUj3b3gzRvwox
T8dphjxruHCBuPgWwYpV33Dy6up9Kr5ZUKkjOta9IuL2qGOKHigU5hwNDXAunS8O
JHYXShTkEndF1XZ8J7qubK52qw8rnqvEGDUGqibR0OmUDgY1O5Whwk6E8ZSJp+kL
s9m0Vh8cbh7LqzOMOkGFIe+Uawmr4z1VAwTyHpuJ0Io3m8BYy+j/4EZGTuJcP3Zj
o229fhjZiLXjBBENrcB55K81q5f0On9EBpFHohSZTNZCDT5ZZH6GwOEbTS+e0Hrl
G2ikPwEqLTKen+nWn/1hQbnvTA+lOPYAO/gb4SR69qJO4/EYJqaaXOTItPyhEp1d
xoWr/S2GxRLOej9yZzK83LRNkgrFgDS9cBMt7PZmiLEO+S1WPfZUkWfK8jA2kyO/
OM7PQhdcfvdgPQhBTKjBYh0pgbOryDPiKyNgSDf6P4bn8anbk+/YKnb2vrNq8AP8
DWBBW1O719Ww9M8YQbz/J5MIxl5a7MsecjfBFdwigvmwK3I+w7Ib7jvUdyAnfGO5
M3RKkDs5aYdxtk7O4XMktKD99wpVdHt/Z6tdt8LQI26iinUgo3G0+pfMCgsb0KZz
06BWNXS7oVjxnouiaTK2QntRdO1amSn9gQQxzrK6vnfUI4vi5JkAbfHOF0puV1n8
GiRltOeOppbipbemsSQUKlMD8ZP9Q7z47K6rlK+VUX+HUtRn3p7qXeHGrMCZ3iXO
Xr3oyr56oDF4oyj+ydMpPSwb/zplbDrUq4ICaEf79P/uG6W8blsyL7h2Kpx+7xxN
9XefUkKzTiEWGQjdBjQVYbH2FrZ8nssiPE2aYb+TrxKXwF1j7UnIRHztaLRTe0yh
P1GfjBvZYu9qB4STpj5Ykto83LugQZGZ5NWAsIULU5CuKvaibr8UMp8PVfBNGTvg
Up58UOZVR4i5sRfWxDPfszKDvn/Do5ljq+cwD5zFSQ89+BzYVqXwTdkJ+y1WAO4i
oEAG5tKMvnuLXZperIrl06NenoiOhtgUNhU6bF9519r3ackZ0fMdp+rbH11pQP75
FZ25NEdp7RNnZAdvHsc6Izo1Vxdx5loQt7PWEXOhwKe6jyizW6u2WPBTwV7Jg0iV
PB05MZKNItxndT7NZFeQCtfvV+diUZDZQhdo7dconW1dLw5IRKpZ6v7BllpYefWd
kdvPRYz8SFZwKyZDUmZgUaYODYM9VtpyJ0JQ8Gr35EhEw0qVli/1Da0hFOGHjNcQ
djmJBNRhK2gP0QvNFkUCPcn6qQfOeklqbTqBs44DxpznvbThJYL6vF6FS6MM28Jl
FGxuss0Vai0j/zA8ypuW/Ku04VCPcyPnaxJ8Pd2CcS1lPpdYY5UT0qtB1dFjcVbP
IrBHKPB2SQ8eaxPAyPGyBrHgwdtkYkOW0j5Z6Dvh9c4sJV7NnFd4g+EnbVMq52O2
EJWA+96JCWFLkb0I/wOl+j0JzikSSQGQmdpN28bACpOuG8YufB7HQH1UrDbEzndr
Ku6b7fx9/Xp8Z4Ot3ZrexVdoxxQ9Jg2XiVnbSYOnt8C0NdiMhqIgXYDM3tzMslIr
IwyTf/8qQiCw0o7yBxj53Uykia4gCDHNC/WnFOgOV2J6UH9JkVLTFhCAppRSCfyz
Ct+7xCMCoCmI4FgAlms6gLufrICDc8lgvPq4CznnyEk3dVxJU8D7DHYNIi6h+jzu
yJUfsHa0TgsvM1gNh8VpJJD5/qQ1sbE4u9Rgx5RveZ3yCTEvPY3LZ9afuvMLxnZh
lMQMdxOUgv9cdi/AY5wLXN0ImS3CWvX/GJY9E9DE9iEtDRNYxiubwRHDJ0TV/UuU
py/pK55NPPIFq1GJ5NevmZbH0q00WUCckqmprlCGNRSosoaCBrNbr/1v1SXfDOwT
NWLc7dGqdMX5tjBj8/gVrPiT/RWRlTiMv0J0xfPI00QqLaXDlcTxUwF72bPr8D1G
Wt5DgRDICWEgfX7fY+B6cbC8zr85+YncEn1SRIsx8HPgaDrFj8rL38pXwLhTE4By
7ZrH1lUhDTy+r29U/xcWOTc9lLfy2KpZWU1o+2wse30oI55hX0F/wzTO1dm/x/5d
8SBXKtUubF4PmnQ0AaudlzjQNNU/wKLlA07bw1mBjxaO5L+e/PAis3UkkPD8mVUe
FNBi+g2Pme5v9bnEtW1MkterZ7FWv2WJD9xRjrarO3Aeifc7smGAcMykuVUDOR2L
qmjbUagfTMl9t632Q+O32HlexO576hT1TXXcUXEpJf7UTy0SQXg+njuln0vjcaRS
h4v0FI0k193Nr4B2hvDHevKWIdbkIQw4Uj0lCxMTlZ/upluqP8npYSttZIA1sCFa
Rhc7sGfKjgjBoBAOHS1FktuIb+yzv275t9GkpWb4JdvPs0PYCFvNGAA73SAh/qmc
QwWqOtIg89SWeRtabNIEW/tcYi0wqytUQJre1gnjoZMPukHUb66oN5HQZyPpIsCZ
nPvEjqBXXr22PbHWx1XHdgTcQhxLPkMXOhBE58qitcE+1iOlZN9j2/tClcuWhd3Z
ZUGGdJWeOzm1hmkDWhEf7Z1vSm3+Y+afLLWYB83WQ44CWA2kI3VRMXQ6i0oi1adS
SDNoGSIHfB/Fyf10M80SEUUyWxh5Il2P1Pfma0SoqMOkPBhZMaeH57u61jjnM9O9
c4nnwltdFGjlOkwQ0IT922kSgAZRdkUFW0yGcIA3hgT74k+WBzucGoDzP37G0sme
IIVNcHvQZGGwKmaFetY4YGEgilrGLmeCfeVKeQGl2jJkokSv1QfbyEoEC3tK7wda
J2fZqGcypG+ucZFdF9l9qFzmC8g5nlluj22ESsow+Krn53SMNWWu1Cd1/lM5fFfV
Iq2b19/rGuv3rv3rtiKBUoGmxfqKw7P0q1hxjc3tyapaC6fY3Ipt8LYqcSeZz1Su
I3hBIEuS9Qhr+KOTQyhLivzBbwTJzC+3gCFqgGOgWxYP84ucNgquv3vCpuxM1g6a
H/KfGkolTYTEXeSQMhCjD0sp0HeMrNw/6BXD6VbPDS/PE4hKEgvHQvTh4l6yL/gP
uAVJj6XFaeHqheG4tdoF/V3nxcQRHWwdZ85zmubmjsBUZN5bldY4IGkae4v6NzCO
bCvvNRaPnj3ahqz2N69PXjzADIRpDE8XM/mW/jwyWXudLjoIwLEVB98suLb4NTNk
FoNyTi8rSggKeQwaSdtX+Rwzh+RQguL/re2rQcdAw1KEdMj7t0KnOn3LgSyRVS8p
AKxTIPy83Squ6rD6twcK2sl5Hm5QzXYPoV8k4Ij0zdG9v26Yhso8jgIgUdraZXb5
/3RAkAaEvsiTn0soyFqcyZOOLsRA0OpmE67TCObTVLf9XHxyLRxqx2YMZp5/n2xk
Yry2g5D9FCtWZSC3k1wIP/mi9lhCXYoOlNdkN0URddR1GR8FRhTFET94wh32e31T
SocAhCjhL6+5kI+26Z9H6XNKwm2wzu4HoXCNvPS7ns9Lucg/Q31RAOb9wPETajpw
f563srJsgVtPT6naaghhJyZFgL5N2idAYWOfDxGp/O1Hzymk36sVpH6tT2gHJS4o
Lol7biuQEWU6tmhQ8hu72aIDDltXx9YP8Fe6UBkeJYTSxE9gwDSRZKIoxJw87gGj
SYxY7+A6K9wqCDptlq7Kbw902ej0gbroMwjF6nyrMk7PzXc0aKk+9VMf6VY2LsAk
SLLKGA91rNhbyS/t25u6oYMjmC7rUEwLA08KMs8Rh02AIoucVY7Ozov55gbqqNL4
BTVYXQyY/E3gwvJPx4dXyQxRvhMxj8moYXzwmaCKmK/RVGN7/q5fMMYyHy2LkkSM
fcvf0/iXVvdTPVDs/U33AMbEcd1UpJzfONPsn3rhjtVtflBzQUi3OqwEyLhRpC/z
F3KSvZrAayaSVMuue5Vl3L/Z9MXNMPXJ6kvxVRDFX4WxNdospY/NZhd1++BfkvSf
EKUmekpDGYfYzGqneFB8ozvF4IEhw/DAwZ+sd7pfdOFY+lL0R0JB6uvubP0PE8JG
uYN++3nt1pH2gFI7jdoPL+Tqkx0bc0kAFGTyc3ARH9SH8MOLT1oI5QYXb53rbd+X
jPAxq/7fUwKmuRwpEaZBE6/VrLioe1YDBlyN/cqDyd40cCqj1Vwn1MWkzuY0fj0D
uyCp+HI6i3Aq7mqArOGCIDxeY+KyQExHvG4pX/VUXMtFvgwRlOHDPJRY5ypcrjRa
VoO/5gxRN2TkPWOZTWzRKpb1WwIwx6qlR5fso5AGCxk9BjNCD9LQ1Xc1pzVAc9fP
mo/pH90qbxDa8/lqUHyhBxelrxzKx2SvuOTlOn18HfKtBU1wB7fpvPMPvpIMxDe6
n5JmfxBCWKLJgxg7hZ1BVwj6MUq2nJ7/5iZwYINkurdo043XzPjS/SfvFH+EUHbI
aHmu30RIc/8r2lS72EFeTOADiNioTx8H9SyBBQ+mxO4/9fNAEiWKx3RqkD0LHLGj
ecahEJGiK9aLM3ALSSXCjOf/CJ7r9Z2WR4twk+bGaTYxpn1dqWY6/jPu/+VhfMLG
rueMrleHdF8ZZPOVnXuuXD94y0MHWZXwKHYUaDwvSqXpt+PJN9RAOV2JMSWgA45z
wnqVK4P4g6bS8U63gkpBm/4MOKCIFtdT58lTcZclT8p5XzYqQ9iCePPp5jtFqFFJ
O1YOaCkDrhPQzvHufB9gG9U0PzI+xUV1ZR/AEHY+t3kBtAzuFesPgSKG77ittOXo
k7sy92uNXD6JrNmD/3sst9+Vva/uUuYcovMlj34zfagBWuUdMaJyhLLyMcojnNpN
e6I4+CyGEDYlxu2KuLsJkmHVslZ22Ws95hVoTomX5oS8vLXkL50r8qJ6OFCNd32d
7J0yG0bXts++bFmM2TuCmRiKbZWbWVsmtGAdHcAjIaCCS/aS//JGgPm3IQCHob0V
+xZo6XnVYYN08YdOp/ZjjKgkk7ACwBGdarBfd61AM6QdH7qfP8I9dQzGJH2lEiFk
/hFxaBLzcXJOQk3Ub96lxSF+5Gvq3XFRGCtuBKUPREEfOCkvJ2By7eIqNXSCELxD
sofdiARX/uSe8U1hbGh4mwwF1cPVTbjzLa11b54DHmsbppxybpjBN9tRiMg5O2Oq
0dHX+ekcHuiEcFnXV30MhWKnse0M+OBIvQDMnSBtuAwuacbyqVnGawPTC7kcJ1cO
3a2RRv9sqk8JFHHVvAjlWetklPM5A1DcRBiIVpbRL8wnqTycv6bqIZcLBNOcnBTC
aviCz2DSO9uf+CCPfUor0h89c5XhAAo7lIozjyqo1IFWTHNld9N8Iv5ZO8ezc30z
vNr2AYIOvmlylv+JxSYYogbt9W4I4QpnyNADhz2Da3IQShAB8AIhao3Gt5tOjeZL
Cm9IUs1T49C/4SYebYCiw372CjcB91nVGlw0TKfWWTrSqgX+D0qa9HwLbd2gJ8Gy
1Ng4NiEBT0lfkDr5pDdgMjYeJtnRMYFAEfoeZJ/iV/qAUHGteJICLLu5HodA9cLb
ZTUfRz3NVB21weNCUad2UxtC/KZVFyUanUPu+l7sL53/Cy4A6kp/vkQqKGTYC7FV
bKHal+L6QOOmrap3GLiPcQsuIWZwu1ezyARTn58aEU11+V6IFKEqX4/9t4GfhqsL
VJc4KXr8NXIu/S2hXra6tjYGwEv0h+v+uc9eOKeq338bQAHF/u00FKNgrG0PJAEQ
m/WmUFsWYysHD83lL+oRCb5pOgdBF5Sr6WIs0newiK0tiHva1S/aZ9u6DLD0ec0y
EkX9kju4TbksHycoGh9/Ary1ySriAlG1u75tTU/7jK/Sa0eqFNZz08T1xZAudPAe
SPI+7U7XHclMDqmpKChkVhNwzLuiPeLmayvyfJA12CGIWqb5W/DhQF59PcJxGSCp
o6EpI/d2dy29PVIrdXdfHgd1URGscmk/PISxkbjSi7cMNlpzMvGo/M8MSAk7gK9g
d04DJc3IHXyM7xCVb/tfOvHQRdVapF81ilmTITmHImjzyWO4FB5cy5+p0CPYsogF
RMVvaYpseb9MhAMKwKu5h+byR1ImqT0r/d4PUW1bNhY/nudUTBY/rtxg06wApyh3
TH4Zj+Zj9RHdEGx/I3TA+td1hjMiVdeTXXI3uEc5ygMYccEskFI8JCby0yud/AYn
smqejh59aoeyJl9AUxkpJGkaRBZBzBVYQsggdHVL2y0XIpsPCMub2UftkhPPZEzo
GSkXWfPaWvG9f8enFhEw77lEprZfXmbT/HH4VEPOMrscrot/YR09tvDaiw8EbzWZ
UM5GgQkKVGQhEcOypG4PAMl71LJ4t8h1/g3HTf9s7umYVLPSd88yJ1p034E9Xy2J
DZVAZDM0TuvFGbmPLpECZLfwXGl0nCdwRPBEmlk3jmKfakv9FOBtR7qyQCFQidXR
vX+NaxSmUyDH+IV+/pZBqH3BBlvEHh7jps/+CFNBaHmUq1R5vAHxh1MmKQGph1Qt
vo6kPCrPTUl8UoqIvI8l20rCTusWXXLPW/1Kpm62QITJcwRDJ2Mfcf7VQdQawhKD
TrShv8JbCJ5ptyaG/TX00U0g4g0XBX6E8Wqfxnk8My85GscMbujnsQPKMH7yaaoJ
lzWjBAis25iwYq8ziL5MR1K+uC4dCpfhnUbI6E6mLDBeNLJF3IDOKUbC6Kzh2fo1
SyFyhzg/7OfpVVwFcqHyczVYMbb7+/mcVY3GYnANQUdLaX5NO/bMXJsKw3oh3ACh
aab+R/ED2iHr836BtHLZvTZ8jI0ete8emGqxmMGd9sRK/ENSiQWqdgXjpBPv90Ja
5Xsy6qYVZsu9BLy9zB5K6htR7r+IfbU7RIRvVBYn2PnF5zo+7q4WtWhi1ytMWen7
ZsrWFjpGGukTK50gmkDT4a0UYKF1YQacyJgBzJyAY5jUe5/B0O4sxEuPMNHE5v6a
pcEr6kXDHWlczJcvDHjZQiTcFuxSiAenjiQzN/vTzQOkf6zt/ZBCSx7AumEhG5Ri
PdYiYYcqlHyHrjkR3MXRW4g+2A9Z1mExcNUbmWkP/wmDJiHMx7VPb1rPsIIFO4wy
FeK1xLr5D7fcp9R04hKfN9Q7Jh9DRKTqrRCDIxNndKs1mvoBuU+ZQdagu1fAr2Nk
oybGGkl4IzSyfFAVqOEhTP5AIDqAqpmD890O3g5Dd+Vk9JPiXPK9qS7zvhprOsja
ShriDeQUfS1wOA/EWWRiJNhPeZ4yNM2T1BRZL+ye1Cb39PfeFxRhDk/cWwU4SEwv
Fi8xlCwoRjs87oWcvM9Ur5TzI8WnXd/AgSHjjPc3/IngIeb9P5j4pXL7dy6Ve0rN
NSAYH+Xc/YG2uEeW0DS1Lss9Av+r/HIryXKyv4mBhVjVYrWfaohUqfZfW5Zi8Rc6
LvD3SysqtnHLi/1nNMdkhHdkqETKDNuJnlFMIKefx5Cr0l1nuuqG6bpbEura/o1m
f0oAZXr/nRsOGIUOM26GgUY/XFbd+j4APUCj/O1WWZUiZHJsannbfyFmrWG0t3q0
SnS66AqAexnor2Z42aFM+AqEguvozIJvx/gZiHU7LKrI+4E+CBrW9gjOWbAtTZua
wKL91XMUAtgCy0+UKAsbilevpCJBTLKZOgmRvJACcVpC0vXxSyHRNLPBjZHz0y5P
OJXXresgj3fr7PEjpn8M2FmPSTNsrCjJe5beNOAFBwjPvZmC5PDA3rzGNc5v7elq
kruP83E3Ifs9sDye3683LJ07BP9zMVmBtZggn61ERmEZZBdOY6IigTM04SebgWnp
+rE2vX6vesPsqVTdhXwknN2nZqvk/kMkECX8DigQ05O6stmfsdRcAeQz+EAHLHDe
XR98xXUZBXpByUvuQXFZeojKmr9+nOMgG0FLqt18soBaTPZM0dmDtqoqjVeK+IQ1
A6iN5rv9+0huGswZcweM9IT9VBdmnCKrEkP7JQZTWa2mRqCOVJHoNsHO/ToAZQ5W
DWVfnkyU14nDC4DM/L7vFs+/e4ADe2Br/UufRP2vCNVrsWy4FzFY2tiwVbtYIIWr
hBwJNSQLzMiiuL5q7D4rLUBbTiJM+ssX+wL8yUocHJv4ETxy8pTseG4mhppGidsK
09AN+dIdG1u3j/cKib9GmajHgfk/ujQXsrts6LD4dMMWzswypF1EWZm8wE9E4YI1
Euu27mYtQD5Bj6s81axm6StzZpJlXQmyzp/fEB4LGfpQBWKWAWDbNwFE3YuNeIHI
shgBCGoy5e8bjxpmiPXgFidOo5IHBk6EPDWbJpN0Tk+sHQixUxxuYu9VwltEG0x7
AnS5lHZVi9WqaE/zlv6qIS1FUyYggKwvQV4BHKBcCYRS2DBAhrBehOnOuhTXuFua
QGuHKhHIO4R6foBLiEJE6Btj1zkOt0tpYKnrCBoID1FZclVxPKnCf0S0FXO9/lac
CG/emWpE4aXglkOU+jr6I1QTapjYc1+IOZnVIKMzvPdUMeV4XjRVx1ldywR4iKXe
bnJSFIyURqt2+t3O5zIhMH0ouinmTe0omv7NsrKN1BDOpqDgNLUhs5Jei4fOJeLi
bXzKh2FQlLno16TwtFIJMyO1NSTxRp2FripOVTRCufS7QlR5ugtjCpoSS/Ekncy1
TlNTSogvTkJiiziEtiFnjbsILTtdPgm+uoGrB9nN5haEu64BZfHQRrtJ+m1bodsX
lDOFpCxmQ+V7V5Si8xLj3194Dgs6BTFsAQYreD6YT0e4NUT+zJGXLTZAobu3Lm0C
cs3pPnivfBt8SKRMNrTb5/UmM+1n3obIJB58iDLY4WGpt8uo/yHE+0FRbWkPIbBJ
CT1NdwJddPVctsUYvBslgLfFMG0j5RVVi8rkBLchTTxbd3tLW6HB5ob89xO9lfk7
JNY3pNWQGOZoz19PNj5DJ3iSH7tEIXTshEEgpopMY1EgjaLhahoUhPTABiJ0p8vy
DBBoAEJs/pbrClazmpVRq4CxxWmCL31D3J4cE+Q6t02ltPdws170/u1ys4SfXESh
73upX9azZK4M2D/Kq3HTEdDMOAbzUOmZXMCQM6AEAEIGj4lRlnM9Goi/Tcjk91s6
oWJDJ6wuzcAh5AQrmatDjKHLZfPIcgg3+1Wu7qc7mF6C0wW/KFbjBBYV5gyd3VLw
H+lglxhrUvyfEk1sjRq9UtEEaSheQXRRfb5JKoaoABxgF5aOsCYATrFX7T7FFzL4
fHG4S67t9IgAD316oYh5VpicXMvi/u9fgO1pqRYOaO+NAcJy1tooafTz+qiX4bhK
89Eu3FN0ojlc6BeUsyxSaYa/lwp57n5w8t0U7PrjEtUAsdZsh8IgDlMs8U0xWgdv
xTVnsOvltjaFecMxVJNRdvdeDp7O3LaCrd3XDF9r6Qq6+r6fBwAQcesIm2/0LUUF
XXi9CXzGQe6v4GBRLOx9iFl6n5vmctCDeQURXZ8W4g4I225kTIfgKESFpWSQxujx
k397tJjqbucU3L7NUU/Fpo+2PqgkFFL5gM7AqNj0I5x/ngrVnY5HOSdI/yBLVd0b
A4fzxelVUZGdwkjq/tSamw0X/N7VWyag3FLXTKmblPc3H4QEM1FdHV34QVxmp2gc
+YikPnvaViiGxdF8m9r7KoEG0oX8cLC+9wXLElvk177KtB7TGiUvhDEpuMqr/7Mg
Hn/pK17YDnBzt1djVK6QXxkgTynQ8gXrpt8u3KouYbcWArDdvillGhDHVBfoSnzw
uugF+0AVf0460qBaqah12YAk8hFsms9hO5lpAzP23enjwm/hlT/VppM9gJ1wdFd7
CWDRw00JKu+JWV49O3dz5O4oNw1BPsR+e5ZtuI3Ma3UiBk9Ti3Y8HZrO7D1YCB4V
0NKZdCkXqHQI3vfY24sZ7qlHRN1McPDMQDO/YeIKlUU3xLPRWljzWRzH9OmPtOGp
404qOoogIfCT5LEsf9B9fsAtWTVZ3zaUaVT6bc6nqGWS+wb/NtRg9UblKg6LfaAw
k1QnxiJTT8NC6jB97WdWHSVSvMqTV4jhmgGuszYjWX880bPmTUhPrehc9Q2TtlGd
heNTA5s/4lJWx7Cm6mW2I4bUBaVoaz08ZCRhPhAYKY5SoRb/mpOSzUqZpJBH0QJZ
bfFXk7XE/GDk9dK1wGFMy+MhviJA/QablYble5l8JUFGfi77pTuemobgU2q73d86
zkwgGAP7jsihuPzN1h0B62qO90pDG2djs+vKaHbVJWdgWsgBCejrdpPNAp3ulf5z
JmjNEMgyhO8zJ7hjt7rS1aje0YVZg+KApsVDBeSvZkX4FoM/FPUh+tTEq0VNKcTw
MQ52Jc/bYVOFkWwdEFZE8bPyKhsjDjMURjmIMOvjVE4bsYEpJoqk4Z/Wp4ulWeEr
meev0E92o1nqBDKjw1Y5rBi85DU3WsT8oAwcWnsOUNcKcNNZQKgR3/NqYT5nsVZa
s9BjK3yfwKHifaL/LQaJ4SnVcmUsiQ53BiBOmBmS1Jf27p+zBGqhdn/ddck/DB4v
xebNIFqGI+edjh1YGgcW46t/qgxSuHzhrTGoB6EkqNzqdTxRdxFppLsl+50xBKLF
D1F1hHL7m0h97A9gYuwc0xKs1Vxc2SQtO9G5d/S65DN35eY9MsH5uBOFn0fEMDf4
1UKu+PtRrMIPvQmS95XWConZmLx67ezs2d/Fpi2/YJrMzZgteD4tHJ1Sen5dWXwv
uUyfNRMdsmVkUTVs2wHIUw5gKEBkaN207hkhWAZkgJw3A+vV4mmCxuCGVenPt+GL
HCFwq5hBZETewBxh5FZ3ue7ql4YdEEEBbQT/Ir8RRj3dTTib5u43ndyI4KRMXQIc
6L46s1QwI1sao5SdpyXquZ521rBywNq2ZOMPtOV3gQuNktjsSQMQG6ohJl2PwlJD
qogI5ZwzXuhVxzHissFHaEX421r9xI8JTOqy4gLzoxXZB/JxD8m8VSmZXoA76v/B
V36H8K3Yf100Xx9w4wBXEvWY8Nrvul53VWiKU9RQcQ+dCCtgbQ/2js1gPX4fV5LS
`pragma protect end_protected

`endif // `ifndef _VF_AXI_HNDLR_SV_


