//----------------------------------------------------------------------
/**
 * @file vf_axi_mstr.sv
 * @brief Defines VF AXI master class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_MSTR_SV_
`define _VF_AXI_MSTR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
TntnlKVgaF5Ce1yagZyW+Z1hVimtJkVp8lZch230hAiNqjQ7LRCb84ibWb19aFvf
f0RoQKUtcStM8jS6W8gskLShM/scksFlErB3hxNqHH2u+FAXkH570D8StBbet7bA
l5EhAIjax+5ZxQoeB+Is4NH+v7CmrG0NjYSk8hQwMjHdpZSOoJXaw4CUU9NmVOZF
pAFnGkp7j9P3DXV4k24dc3tvb3MJYY9JfV+hJ5VXyhmwozXOrk6hGladUjYBhJr9
yRPPBS4NBKs/JpHSyEsKrpHEGDSVuNyuAJv/+RbVV7dYDExAk43EOwglaX6UP8UI
g8P/RN8D9lqO6XS3bUU/QA==
`pragma protect data_block
dGOqZF0zQXxXL01TaFf6Mv6ud/XZM9P31/ghzezjcBRx7Y/IrBGq63MtZAZlvJri
z+mdKIh6BilsMdriWxROhQdRIbX+FjGSURytpcBORCviScWAUwpCdYh3A9R1YPF2
z/DYrY8s9jV0/ZcD0Id3nsNNM4LVi33i1lGRIyyOxUgPkA21r/dqj21NpvZ0yvrf
iXzxMWOzS6Qtlw6J2F4Xx7Fl+yllZTpMZ8yMrQkF/RrYRZq7kGKHML1u52lxZKhw
eIj2vWynXSZc9Nrbn0mQLwexcEN/utpUUBBXkzGz1B+3zFb5K1ppZWqdKSiAEnMM
UtJ24fWCDlpQgOHDdvFq/9Q2083mX7KcIFdgoEioOrVZfrni3KWqo1iz6kscbSKk
J1jrPiwaVWiX9Uo8UYvYb3IgRN33vw0GG/2ltSWKj6izwESukLU9W0NrRZauSY4E
7al1lFVlXMYyqafOsT7HSAF2FF9aehP8sXIlijgPWhYTiJ7TUUp05kmOh60CzDaV
edBD5RaZeyKJnCv8rnP+4e//kZNAht8lY7uRnpZJZ/vNmZLjg5YnRDUw0kxkTY2h
+wlxPWfK/ry2XCJ0Gx4coJlbVSFvYK6DhyxSF0hMq6fouT90pZpOhA/2MVC2Dvvy
zlJba5yKSAShzKtJakv14W0SjVqL2IFoC8k3Z5iHIWqDCQr9qwEnSqkRUf1tUdEm
f70knWVBZUqWA2wYQkU7iFjMjpZCsPcJ1PlpvxE1fKISyldEPuTTFLupUEOUa2k5
gEU0Gmz4Hufy3vioTiCn4HqYAf0zMJ9mcnn310p2SsTE2Nk64fRvG4RTExeSf/Zs
tj4MaS38BeL3NyA8CGdhEmFJWfHf9Tbnqbo5hJH2zOL5vkZba48K8UJ3Y4dfCVuE
mGQSiLkFFGxH2/QAGdmYuGUZ9Ba5hJG2b/yLrSKerDO7vwn6nm0CS5R8pljxJYaj
ntK8LKRvwVVfNVl9usuL7ZV2of8P2CqmShXqWMLNGT19iOV0O/4uPbL4F9m6fkCn
swPfTtGnzxP+qYsyeDDydR1xsfYbIw53tNMjiKQDjmchpi1NwbNgBNHAa+sf237N
O8BDgFv3K1RPCmJyEwjsHWR1yRNH9JfzJp/Uh2k7eJqW9PzjCMqhWqvV8bZp8vkh
vUOqZmazjI+J7pwHURLJ9GeOjFZIzl6l2w+TsMu74wskYlQ6D5kc+rMJ2tD3DB0q
KcTzkhfFDlTNPBeqKmdFFVKuzPHUBeDA0Osie8OWUJSy73zL72pxZD61xsl3rlpf
OTY9k3120tHlO4I3VujemgUUS688u64H9eTeOUHVDzEHaFSJbLwSbqShqzV8NioF
L/9OUMmRuhtT1WDOZRbyXXXPqoQ0d617VC9Ky8OaHfhVY4dXfZMTHT8TbEQEINaC
aplLy5CAsLQRKD+MkIljDKQj5GtrD9VH6Yo9/8EAGhu7PC2mQ+bgFyLj9eJU5FD7
Tqt43jD0G1/dFutpXUIBFyi1eEtzqJjSr+Uo+hcF6bQ4T92vmyHLT9vmHyv1L8g3
JlJ3WJK4Jtnd2S/8+k10UPoQfA4wzv2hIwn6jYHTpNEvtEUUGPO2NwG/4okko4up
pm233d3oRigphkfHWt4hbeXlC2+8AAdq6hX4HcJQwQw22wD198IOTPKCSgI7jN7J
CCpW7akV6nTZKks5hoB5KkVEc7jOjpo2iG3LuiVCaG8covU6a3lOxdurnhdS0tdT
28bPNTeOWib6ggYizONScqJsfth19lwnDOWe+DZVkrC6W74nAAVFqcbVgY+xDv/7
OOLAoxOXuZCCzfmYueejpxzB4+yJ47vmMlafXPYA4Ev1xHIXrLrya5TJoLDhpfVk
2ml8qQHkF7d8JgWEYkyUlns3NtxawivdLZLB5u76R6Eid0ZkvpcxK0Pti90Q21V6
9FqFi0+BUUwZrtPuy0QDfFlcCAqtc96i6cQBdv36zi0E567ru/wChB2FPUGMAnAg
Km7o5gb4cPwPiQYo5rio+mReu1ZdI7bm8WJaIrnhGeowcM0atsnvoasrcuc0WLWE
ZX1hp3MRNmaPgoZ37PfcTJJftRucOB2XOJ2DRoPnrlPDKlPSdXw24toIciuCIKWM
MmTyurSSsHPhsA/HWu7VfhAImprDSq0I7z2jd0Y7ZxzphqlL7C9W4uT91/31MJVD
nvqxSEsS+kXg359haZdL3AT5VLXvzuL4/ni5dR0d+WWxnzZBmfxk1/b/3oTOLsZD
RuHH7kXos7Addf2oM+cIdKPnVP7eCiBTua0Q1w1w/iN69Trrtw65sGavaHMS/1+4
6wxczCarzOpg8YSa8f2e/JdePvS/UAzFsuL2PwFhZilrtwZpNH+MJiGJY0IRqvKM
TTvM2iH2lmjl7g5fTsBaABaMWqnX6nASz2MqMCUUf5tznNP+CvbiKx/2qLUoddJw
0mY83cLdEQ1CdakpU0BgPNAV2g7pqlmpybU1gtcMnu2TZojeLgRWkTehAx1Gk2gE
3nvuyyu4cUweRxiNG2naMp2qx1hJgij4MJDj1Vt51RyqR59ONFaxsr7ehc///oqG
C9S/6PBWlC5BGvOpx812xYdvdDpWWnXK9OcfeW9vAdv6FRff0p2dAQMrsVa/Anmd
gf+4R3I7ppoPeuRazwMFtQcRSGQwe2phMgKAh7potsdXEqiIj5BD6j4o37gJFtwC
rXMJoBV1PQYbK5eh8krFaMm13bBnCRxiC+RErQTP5rZkhzaNtQPUiNOl6dZ3msCO
9wK/waYjoSuzWMbQS0v5n0ahDbV/RB5WqIhz4LtCCtDkTmOQjYmrR/9KFAiR22YJ
4WdYTqkIzqzeRKEeuzYGi82YqYNs3EZQJGxgkFS4LgTdrUpA7VzgjN9BJk2KRpUD
9T/99cGnz23YwhiwiCNI5l1oLO7Mcl+4pUAa1Zl3+OxO6AJcywvIlhjk+lnobelN
jojTeUh0eFUfuJdSpyk5Y8DrPzF92TRhZtWoRe+AtryvJ2VzngfwxQvcz/qEd3Ou
h1lfe25EXvhJkR/73PMyJ5t/lG73j61lfJBW0EevngFRx/6Q/VxmRw1fuVf9KOJG
x7iTCK5tNf9aO7gOcVauCmCVKwAKEh/LVTf2c13vZaDbe5vH01JHlpCDcbHuymjk
1Kifttib/ZD1dCIcFE4Hcv4NnPfPUYcWvDwaGJMKlUtIyOlFzZJiRLPKg43TFWpr
ISzbMeQTmncjpkMO7q35MPlIikd0dIwFiMVVqQoxKhkOs7v11WfsFEwRDnL0Mu57
VXzbc2QvqH2LntFuldjrJFGiXYS61OIv2x8y0s4bAeRMdNEe77xLpSk5Osc4mnNO
uDeQDLtiJrxSvis/zLyWdBkbbDaLFmdvfp444WzILj9y4B/oNJiUCqiDU5QBy6jK
pzqlShFba442HG3aIuXTN8HO3NCqQkJAsLHSb3qNx1/uuTKWmmSJ+vPXJaeUXbS7
TA0QiIQQ3uv0ExePDrDFTOYpDnjm8cUAVdOHJ683LOHcnsQotkUT2+B8ziJc6GZk
YXPl2noUrzM9HRr0eIS7MaMehxixtd8+DzIFcaSLR3ViAFlSx5m3YUe+thLDC8wk
rqbJzJZbNhNFKOF1aDfs1itIArZnwXWmDAz2zMqCRcj+lWAhKjbczQghq6dLfWag
UIXb2vfHjHR3q+nAeUfOVDF88Yp+Gwzhg5E/liLsAHeApUb4mfZnOleAbKvJTg92
ZGiSRRDW0SDmuqtpQWMQSi+tA/yv41dTz+PqpAS6Abo6Tgu04KTy5j/WbghqVXkA
sTdmZJ5Q4giAl4jNN6m55X2DRGSAyIarq2kWJRZ9UM9FW23dFBDdkLzcBTfJi2GF
p2oQ9OA4EtNKOXEg9+0nl16krUY8VtbdnXipXDUSEKI/r0UM+4u7ZJgUd6UwNfJt
grzgAweGvPKsIqlYb1jhy7p95BsmDjX2irEhQ8ZlCowkaUjHCH27zgO9IERLOu7E
lJ1x/42visuC/huuuKrP0JMK1oTVbHccgXalMAVkzZ1B0ANyx4QAu4tm+g0RWmBO
8ryfPuRnB6DWkzsMZtmRxsEyDJj6vNyuUyDdAOlF/xDTpbGqxnOPRnOai8ypopnq
adhZplxfvWgap8W/4xf7ilGlYVNlJd2mvTkrC8kRSE+eLmYBX2IjvQzqJxhpLSB+
ldEO04Lf23I9rjAKb5Mj/ivKJkOg2B/riSzA6DX2mubpENn6CSdnEkhJOSR9u7SH
l623o9DE5Idz0LmVH4K605/g0yEFh2Ke5AD89e7S96CeAd14CIp1XvayN/M2R3/y
XQqIVypaQVbhBhnhDHaY8Rzknw4mm25PLvQ88+buBM7noGHYFhedUVMbSOxdiFdk
9KnmpXoN7cx/bo9ejFkfsWnu+KeTz0xzbmkvims3bAa9wVhmjth+S/JDMi0mwV4m
egbulWalb4Yg86MgkgXtGV3QoJol+tUmdJ7AOLnyFw4PHK4sx8AIN0s/4iHqbgLU
c3Z1LvUYP70hLVKgegoXblOHuCMtU2I20ux6BLa4ZsnJo9IJF1T8egfp/zn0ce3q
7d6plNezy8CEW7PaPqxBbPOkH+tXnHFTVQVJmxFjlBVIzU6LZYLFol+V6/yZBy3E
QQd5mZHEbTrAacqblZqGAWQjwfnSfq29UgsV70M/e0QHq700rSiRpED7ju//YV9t
ER3v8FyU1QFsVTfvjpAsxJoyDtm1cQJVMW5Ev8WXE3ABYWxGTesDE5PGRAUQOLyE
9O6mIz2+oeGLA1twl/xUodvN9Ffm+R1n9NoKkrO4S4cTwes75rzTPh4bMxE+lCxo
yaSkJwn2dKb5WeTA5dqVSR6XIyJ3GW5ow2ksx24QrScVhI0UEwLb9LnfguGdS41B
K6EbZMlN/hcix95a8iezPVRu44L5hKUMAaMYyw82d1OmQRB7dTepsVoD3iBn6Qoc
LLE6sj6d1J7DQBStkL7BC1PGrH+1Pc4jWp3obZ4pvogcd6bI+BtbqASJ0i8YeLYW
A3LWG87GZwOLQMZuKO2SFbG4kRYB/7Ik+HlLT1kAT0YOshBylQy1/+Y91AdLmp6c
S6vWDFrT9sdVKrzH1Ia4Q5cFK+4TLQcuNKcdCJook3pkLL/benooToKum3ArVMmL
3PLQIYIQ4pImWaPrGn2goQzAqy3R/4PR5eMe8qKSpLGAt39xMQipPPBxgo7bx88l
xgd8D/B8CcmIqogswN/7yJRGXyUJ6761En41Cy+Ihyd9dtLaWA732jJp7/3FOVRB
HtF+fIiHVkQT3HzNAT3onlITO8hzDg7rBQ7hxO+SluJGC4HhtizsUIeDFf4b6t8U
fPKaNQW1/b5Ku/C8tcf/vXj1Br+FSUA0UiR1Qmj4NqnGP3J4ZpePulgWXYNg2qnS
ReyaO7l3yqAhpUbjErbl4gvKTcrEcD21tQE+8u3ByG+hpaKDHvUjjvW/b6DQvHXG
GhhhaOJUkCXxDTY1Alaq/mIqQJ1ltjri2ftRO4cl6RxxFIythcslzF/A/m1CVUau
C1ksZvHaG+Oyb8pDDTlxP7YBqiQgsnCqSO2mzjgLh/dNDNBlTq803PRd6RUlJ2wu
IYswxPSnTvSQVObhzTIlnzaEgKqUFxsKAal1GLLIsele0iQBqkKtf0gefRsE9olU
8hkakq9cPXPkdIezqYBa36a/4B0rBoi1P+wSNRoAVxARIIT3YmgKtTwA1lRtfZN1
1e5Fr5UhnE9rTPLO7XL8YMPAkIaIH0Eqjli14tWANtW+MQz+dd75xBZcfnsKQlMi
fAJjwuLqXtaIIR4WBGi+8QUa0hlt2D89/j+pZ5E4bilNV+ME9Faezt9C81TJ4/m7
Rp1/ldXhNvH0QE0xp57WGbTcx5iMlY+LdfvhFQhteDCaE+nbG450BMJdVcxM7TZs
H4gU0Q6dNQO02Eo2yI4LMFhI4YLaRC2Nyq2eN3jbsn1jBVXZ8w1uvO4mMhh8zzH6
GPV+lJUuc+U4nJx9NSwV1YZXiKJFPZximX2kpCapjCwUCbJkerUeGffkFi2QQH00
tdJVVmVgwaRpFdGN+uQZ9RRXeHmDSd919Tj7PSblSL3dT1/i6SHJNT7mhyxESjlb
70UtNWWx7UmYbWvE2aODT/dUc34y6/KsqYPqFNc8ltLcUDfxUqpqe5vkNWDMatGa
ip/iD+B+LMWFMmWHrHmDbSi+pOayJ6v+wEwru8hHyHUb0CVBCJP+3W+KptDLvcmC
AtcYhfQ+t2BlUzOwDTIgHlHCSWn6VXpFo+cAOuXFj24aH01uyzppHYd+a9eS7PRJ
CHseqEwCViwJiS8jBRkKwjilDCC/HCHJpfBh354XLGMHAdNB4AnBsXNbdqpdAqFz
lWAeHd7oooUVub1L+wDSN3gD9GUIBAAFKwMhheWeApB+pr3tRn+4id03sWwybXDo
quZx+I/07FCH344lWCPsmeFuNfBt4E/tC6XIXnnpMaeqhJzgevMbQA0HB4Ex9oMV
qSjvPxhNSXvleslmw9VJvKh94ZgzrweqP95aLmIFwxTit0f5RFAPWkxmCpkLTmfm
dmDuTpdRvZGh+TWCoLTVRSpW+oKJgmbY7rcptoO3P01aqx0SfF8icxOWf49Txo7q
dQhxHWwzFHYr6PURMUgZIthZ1ou2gXgdfwGgGkMeiyYu8NUO7qvUuSSXngX+KlB9
dn9rTi4wkPFJLQ+w1NTpQocZtBMicxi36Ofh1cZb6sUgiHpzP8wLirRdSwefiYOs
sZElT46/o/4ckcxPAjc7GMXealzbUgkM0OeHo7RC224Uzj5QF7P89HujYM9ZNKIx
RBUrNcbhDEHtf+WfUXfPK3he1LNpotKcfx2kz61gohp4bAQAOKT/hA17fl7mebyR
uublisgowtBhLc/NsoPt4WRbZ/5zOYCRIta65i1Pi9zcTExpZXfHo583QWjL13gU
VSClxEo/hQb8JcQ0xS+D/wgwYsKRDE8cm7IphXaWgknR1sL7bYD1DSFMyR0h9NXy
RA/Sjwoli1yYYnzqNoWfrssyEBJWiQgl/DZIHKFwXNFU7cP5ttBsg6ZFlgmUftfF
zeuxi2zTv6NRpfo2goA5X/qKTAhdM+VBOvKXCnd0bI5Eqx7e2eLh/fYVmgY50oL4
L1dkSH9SpNau3sXJUsFGL+QJSMXCgU8+WkOgp5ZpmIU34P2i0ffIfZ/8ZnWqomcG
xDspkg1iNWKQkze4Ir7Kyp6pfS1tKR7HOOOawB5s0el8vv+7M0J+fZmD+E3RF1js
Nmwq38+Cq+wAcQFQHGKs0dfRN9G+/J1Y8jNuYyOnwQDtoM2CoPpowE4NmXynWrFX
+v8h5xmwOQFZG246uxwQ+7pgcXXGhCWiFHuYhRdAXpfd3GcsxbF/UqWgFsDBdE05
8+OVOm3Z7f+bn5zUJGPCq9pEcjQkHJsBJK0dZlByvoypo9eE+dv1HAIjzDS5yFtL
wYuQAw0UJqC30d0Liv+ffn7zpajZJWQb2CsSDERFZAx40Vb4BJLgbSpTQP2/JGKy
7fz3Qc40pFbELkekbIr51MxkbJD9OC38j9QDn1OCN+5yBeXWH9SWjJ6UW5ICyu+V
wKWgZj09nHDtD+1xQ9c8iwgDjYhjVJuSccmuPbJv0DSDELR+Np9oxrPEy6kCk2LP
fms9vg4RqUurMyNynzUlNoYqlHC4dB6VWX55a8gCqIYibXOYaguGt0BeVDd/ugOg
i9cZQHzPzFdF+n4s66Ys4NZLp7kHqmD47eYLLpK5gvMjlDpip09WbDY4v3lL15A2
gDzp6mDIeoxPH1s1ujCciAcgkBAmFmc3OVXw8sLD0p5Hc0qeTnXNvsZmIq4dr7sG
bvsK8rbCNO8Zgdf0110Y1WbZzRVoR52f/1aMbLMC9mgYLzR3IKWOW0yCxW9KIr8V
3N1yN090BfGhFCEQ1lsjj7OuimAAcrizuKsbN8QuoHUy2kChbH0S2v6JggJX9edc
EPgoJWyjWUKjCaYQeubmp9okDpT3MNCScWgaxSXzbJDdCDyr0ggUta8VruMDmVUm
3KDnjiLJelKoHtPOFyVowF96aI0Ylz6YBiy86PGDmnAMMCpdFYyWCX0tVOxzuX5e
a29Xsu0R2VSmrxfFNNS/5+ZhWnk6c7oealCQaDmHgcA54KvXaO0Una5RBzmN/hwf
IPBYZBnAzBHrQRwAqDStqyQYWTYcT8UrAXcM25pnVhINc6OeBnpLjihc6nkCk6f7
/dMhofOO1f3TZReBECseVl1imKkQOgXlDqOzH3hz3UKMIzl78zjumPlM+tW5mCvo
JOEIVUzZGK0nO/twXrOiDTC68TDt4jG0Bfg+wNZzBUbcBhtpbbtshAn49vddkxtL
mumihduNhmCTDogR1bif0wYiQUYmz1kOXC48EFeC5cDE98NLIJDTXVIAMFHkiWgR
eBfWpX2ut2Xk9Gaqsra2tHvyC/e7aTCCM2PYlhiozfHFl/Qao8lCc1phLvkNrzEN
6/+y0nffFDEFBSXEJ4Em6zAJyTPUMuFR8vhLJHFtvGuV0Gdxa3G8Ae2WfvI6XEfq
e72edmWePPhZbhyPs7nziaksP35kOg6I3ALooiLgZ0Hv7doLqyve4WEiXxVw8tHQ
krkmg9l5QCYFwCw8ndOK4duw9SI+guFpdbsguc4gR/UDyRkbX0qufnfH7YZvf/AG
5WcVz46RNwCwOfJ6ZLUbgjPcwZ/JVwp1Zzfbvgssa7OlzyEFn3b+6dD2Us7ylh0J
N5ZjiLL/a73UPIZDXeX497JCqNrstB5cjcqlAETSYUSPTMIdnrH0+4fGmZfrqVBc
Rjy447A6Zvt5kIGrsl1kvKrWqSXgTM7JgkEpunRoWxvZc6iHT3ywIVXFnofgLEMt
8c+lDRorKu/InYVDLDC+kyLJ1dKnm/2Uex2733bGJhDI7u+g8dp3q+tkwwKv8P4R
g26TyP10MZaJWR/Je1cFzWrbBF9jNW/12X1KpbJ6upECHBAmi1Sdbb/KCc7N1Ev9
aMwSEhXMYh4ncj9O8Lv6ArpetZAHSo3Asjoz5lB5u5WsYmUXNpuAsjEub4JStu7u
8mh4syCoYdnAySvh8q4KDkrtkdbCrPBZGPkWqPKJtz+T4OlpI9ExcelY9pMKYsjX
+nsuQ1+Y8J4bA9ySDzhiANtf7uxYmdrLbZ05W9ar1BWd38dbRb82YOtvl0eKfNIx
wQfkdPibXtUmULtiKuPZKStSbajfma1rvIgVR3BmisdWtkEE8YpErh45AQKNwgSR
kkpn7Sxc1/VACr4ZeAmDXbeFkRRnpVuWoTtsRloWevStwwFpdH4HuyLGgow8quWN
KlJdoRJVSbazqZKiWdC2L7nwWLvInScvH9BjtgslBpwF04whbnfc38f4dVKlCjDA
0A3JtKwS0DCwkajGaX5KBHRGiOXFvfdFKhVs1hzkYk37U/zqoylyPx185R6pPYXY
qZZnvXtaiWvbz3EcaE6V35TbT07vd5Co3Rth6a8/W3LCy/HdJLjP7hLQ9skT1NZ6
2NFXEbMvItxb3e8e5bCSYROLdZ41c2gh8WYEEY+3pN2tFir1wb0esT0osENmb9kY
bqde82/Zv+X+0VAgqtdQ7DhzaLzI9ZeIyBCNVb/hVShDBZ26PvmPp6ZrFBj14bvH
i++sQsaitb/hQZ087KU4N+EW7CEJJ/pbnoYwyuKaJfKVwXe7ki9hm18wBAcdiAL8
zxrDtHtNCGp7VDtYspghnXA99t96nWA1xDWlH2ob4cRaFfN1cy9hY39gleXNMyh5
n4Nof7bXRsmNgCSx7ppzITcIalCmEXwyBwIVsj5PLdnCC8w1jpD6AtHx739/jnMa
FCa5C/ptOOmSZpakpLR1nid0AaqXNV6snmS+8Npuy0vsLUSN0w2gAtska/KMChbF
lwVqmdTGDH89hrAzkBb0G/NE+jXoZ49/htZq5xv5y8aogAG76hA0Vm6/ZljxsBkh
5y/vFBSEd6KMw44kcMQ25xcxjsMiqT3RNmAMTilxmi0Mu3+zqYUMfBE6aeHSxPWR
MR4Wc1iURHfegZg2EqdMgnvmRJuRvKy3t7pJlKe7DAcbvbDgudm1t61JqDbIPkL3
rnPQYFBfYBHfg5vjZ4okHNU3RriV2loQdS//42y6J2W/FA7FH8hOix0n6IDj0DDo
VUMweivueVmsKb+PvJye4DoD0AeAqf/VkJYUwCrxztxA1lss9HuTYvjhIru+YNhj
2iu13h3LtS4q/xgPRjbYMn4u5ikrC7eC8Pze8yZbVn12HU2FmTtJgK8uqAz9ztjT
h06GaEfaTV9rb9RA34E2ZOZ4oKJn1fTur4FJqoWC50iCxNv7/CLuubEJGNxWvGUy
GcN1RSThHrx2J7pq9sPX94etJC2xgpqB0zfgyOoYr38HgkN/BWReQgPzLwZrc/yB
DyBJKZdHlIWUBZruaL3Grq4k2AsSda4MVE9NUMykfTM65pr4+9auhq9yCCVfKosQ
pvhiKol5Cyk1Geh/1Q2chpe/lpqfmvy6uxAsvJpy/d3Sz0YrxqF1eN4cObyD7EA1
WnrLrcycYYAWiRK5H1nFbUUARBS6P6WNc8osxfzLmimgrTngJwbjQHDPNyevSTwf
/Lols1KYv77JOa0q+Dj9NX7WN5FhWsdi4ycw8VoYNBliSBt6IjRysuCyV+I/wNpO
j1pIHQCv0QXj1RtxjSl3OGNCsm4/ERFJBXxacJj+p/0dpPNpr9vdowHukv1DIlbh
rOyDyfetl7TEPggwzshusD+vamIvl0DKcuYFTyj8yKvzX+6emeVVMSRkG2rYxUOW
I5jN+Pyw+PBphXsyGQVfNj/pNb/sSBGHBiJf2puGEj5Qk9hvaLF627reSUWap6Xb
AtgQiWLvTZXsLXUsZwswFI5spfrLQws02RJ+IA8MdUMxqFYoVpYEhPvfOH2IS9FD
4rBo60FDK3/QhPz5QFC4pzkbRaecOtEWzVr+qww0SR0Ow1V5GpHil0UD39OClL1m
A+yH+jNP+5/lngERSvzMycP3UepmVIDKe7zUYb11Cq+KBujZ86htlCKqq0OgR3XK
2GwSmHK+4/V5YOe4rdNUWPgTv4kKJJm+6iMehn+UEEchVXTh/8y1Yha20Y280Fp2
VlsywsTKgoLSHVvZ5aFscHqcoY0bULY5NSnKzC4JFH2uEVgQb7jPRG/q37MiZktr
jwdPnocuI1+kJPhaNG4fVhmV1VJlvfO5oFo46qY5+YWFUW3oWHIg4YWPT2347IP0
8c5BgtgwzO/YYIJcUZRjyFbxsQw0x2Qf3wzGj/woeU3GizDj6AuWVFW+MVF4Ud0D
lhGYr3XAWk55cTylziEVCw89pwxu6iQDD5G28yaHOrSP3LPzXHzwpMEM6ws2oF7B
lLsTe3+DDYi09MQpDNlw7pfeccBzYyRNRaxZUVQ4Ags1jmu9XySj49FBzyQKaKcb
JfkBFEU7q6vbt0SqgwVX76tP6wSCagsXxlZOlAFkcrdYWkgHA/YZtuFk1uFEproK
wGSw5lhpcYc5DWuInCB9G7ZB4UGMOhHPElif44XoSZobwGN9t61XpEklWpCWEtgQ
HQsXrCVDoJEcEg0BQi4UrONHUYLfsNmzhNqrePgL5UWxai0bzPP5zvxotiLkhHdq
I+jcgb8LVSk4vIe48SQFsAcDlxENIEINQ4o0+BdkK8h57R5Kd/t8DHMbY3y+CcZr
zAseE3Me6084/atbm2ijj8sxsQPsewGxGmwe+oO3B5lSdc+o8pW+awO3DgnnwXqC
5AeZA202gaLoFMJJa2TS+89pQnj2RnboT2d/KZJkajJR5KJr3mUNEfD5JbzVHV1+
Gpw+5rlY4r0DhmmLegBjUwYCJLvHv/I/glwzN0xgnUNAyYkFisX8wy+aGAHKK2d8
r9HXuL9054kr5sJvcSacfl44mt46cNt5UzXT9Pvc1dIFJmcKIhOSQyoDsbT5mSSB
7dbh3WR/u5sYDK1W63k/nRAUIaunzlH9/ggeGUlKV5u1Ej9jRrWIEdo9X1tgpO7u
OwICY1unWg6isG7WGtcteBPrvARf2bTLYdNh6eZ1uB1kfu+72D84AbgfbXc7Flst
BnTZjMjoes1scLGybB7iAvhhE0OoAJnHZ+g6yrMDKqGgXPLgmU24jFdeaW7kG7W5
oDQ7whDm7E35evMKkb8pDkvF6d9L/HmppxCNJvaOQmmmTlvcbXiJawiH0H3NxMI3
V1CZ45xALrvnLCbZde4Few==
`pragma protect end_protected

`endif // `ifndef _VF_AXI_MSTR_SV_


