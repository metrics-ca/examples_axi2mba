//----------------------------------------------------------------------
/**
 * @file vf_axi_mstr_hndlr.sv
 * @brief Defines VF AXI master interface handler class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_MSTR_HNDLR_SV_
`define _VF_AXI_MSTR_HNDLR_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
EyQnJHmx2z9DD18gpCBU2OZ2ZElsBoLXZmkb2qgQ8qMPv/nRkiqdSsWeVda+/QIz
yCNI+sOgpUuRNpVepg9rh5NetmzHJSZ1h5NZzRt2IfncS0N8MqHjD6uNvqTGGwSy
7LuJPhRQhwt/SIMk8TmYjf1xZ5qz3+26IZhbFHrJLykIvmn+AikHPI09APvAO28G
hTYUbx6NWn0iya1gTaCW14lFblf4zAWDQjIo3t3kTQnR015FFhZJKBTRNOI028Ef
ncksBGjmA2edlmoL6V1wpfbv5mogzjnE66WVud1aAzjjTqD42RNBYmvK32CR5t++
mI/yAKoem1YKgQANLX75xg==
`pragma protect data_block
/3pEKpXGPBPsnEIkGVI8KzDy7nifT1K9oaDPzxDvqsL0iRBsggsLy2EF3Kpwp0fn
leEITIMQObrnGd/9X7LrV/5A09P0uVvMPn17/OsbqrrNhgabHK/Vgo6GEtOZd3ok
zG/1O5VHVVTahf1EPxfEpuilxbZp92MfmEAralALjg77ScUFLaQUJ53Aw5l6S/mm
XSPZAIHNMBQbUKfyOa5/YyHhazUrP8ign6Y8Y7UxsqvPgnEllXTgi93uyruFXthu
kj+OaCGZdAYDN8OkyK3sSn7eNydkjXxPHJPlsN1vqha/hW3CpKb77J+5Wi5DSV7b
+0/cuX7/PsNwiH3LvCSx+ejFSE/FUSSWMHqbYfqMq+3J/ms28fR1OoGJmpdzSVYb
mfM8yF/r+yoJzjAJMP35dqJkQFrS79tSY6CBH+oOk6rQuPc0AoMSRSBNAT54f04z
9RJMQw3+Udt2V7O3qezZNkrD9wmLCMc2N7q/Bk4YZx8SCk7+6PNvAEimXfZtZSLq
/BZlI4fYnZENVmJEehmuaWvi+9rZj/CM2JfrTNMLZkuwmtaqzOaCYwoHb77odphZ
PySFFlNAOg+uNJIVEXoPiQ0NtFfRHheW/cFtFQy6AkTlxlFRORrgGOf/jx3UznSH
edwZrj5zwehCiaHpKC89uYmx20N8BZe7N8UFKb4SaD5e7fTmRE0/tC6wlFovCgFf
9Qvp6Z8/GNXZPtK3rbrqsOUETRtNBluySfaHsQW8gZEoqQMv6dDBlw5aTH2/BJ6K
xyidvVfHGQNFTpM+LuHCDDnYEOTyiYJGhp99LInYW3Ce2QS21uFrI5zKx6DOPRN/
RccYfXPbN9sOE+wGxDyq5BQ6Kl81pdHsdqA2Ryd6I9jejnW8+mQtA9XoENj8OH7R
m6sxg6DUDCt2GBumSXiTQKGQg6Bw94A/ujmcShr92ecXmMmoFvJAVNRo5CBkBI5E
DC8c1w1GY12pdQhkOYD8e5FlGwAgCuTJysmxQW2vRRVMaFg4tIF1eurdItOV8WsH
6OYEIfgVWZN9cJ7d3BIo8NWkyrrvzYlItRpsfcWKGrtCTY33zBgSMo4HFooq/kCK
+z9gSfLQdYyaT4e5ZNY/2fSFgTSM7I/95GTX8jKJUyUIsoxlvyTFGxQyxLlxSeRi
iJEQ1EqQcNQ8wFO8q1k36rU7vluWjIrUFV+E822ZpCtjVvzT23BLB7TsNYBlRh1T
WvA0NNvAeMxz+j4KyKU075bWj3tt4/gKoINxJxYrpkHbdvrHr+DDzW6ruo4Clf8A
yahmKCsiFODgTXWQo4PoU+h68pUdU4TVZnw/bWKeXtPeM9Tm3GOCT62ZLacZ8ltO
enShzDCT7SAWyuk0dGctxTvYD1cZus4zFStsS2pDAnGrlnRh5PxkBaOr2RdYtbte
XyZlyFRe/BeoYcyRLYg4HYsMRVJzpIT5fvLygYrRVtffLems8NyWNmBTDglkVPeY
UKR+DAoUlK9Rts+A0lo1Mg9bFDBpuAkFetGdFxC/uYvDe7kGbMC4r9/aLOpzVvGU
t74HckKboBivqvrYAo8oyhuB3G947sOnDStN56BtjxbMn18XdCM56C9kt3oVMBIL
Hm5hDKrzYN49/g6vGMrVpe6ScgVgn/aMFXVhgbWygcFi7oDC4pZLEz5DAEWh0fgI
tvUn777FsAI15IJsZIOOTWhJobWTdrXJ2QSkISaKMH6KxaAGMFHtqvsogzYi6GIK
S/gQRHgzpsK07vGa6J+ZG1YXF3cyFpphxTuFsP4Ew4L0gUfmIhM4IOzmEXw4yRZI
2epEEMUSbdhe+OpiQT8GWmBCMkh1YATnY7RHyVrA553qp/oKo2/BdTgWAYv2pFH4
uhG/4HBGuZ/IMkJLPvfYPsTAmYnUXu5OJoSypnu9GgpiEk6w2TzgB4t6ksaoW/EV
db8xa9dBHCIsuNMpg9kqMVllIV/90021Zii/S40EuMuatgxn0C9WN/DG5F7xhGHh
IjSWRqzrk0/FJ5g1oEI4vmR8vA//p4GmORnA/d92lt3nlqO9S9nYtjzkU+VHMCeF
LhALbl6Aurin/kMPcb537wfr66kpOcZa4blK470ulM8F6rM7KvskUyPbY6NkzgHS
gRSUVk6ecTqDTuvJ4VCaR1ri0J6ilyY+zUJUVLQgieSeuOgf3MrVHQxIWPtCzv62
l7m5bZhk4HR75WoKYalZ2fCtWRrmfldPhBSQIwHoSI6ZXbM73hWzEpdR8qwWs5FD
8qwAWeAgO+DvpVkYVHis5bOT2Pwgf6adEOnRMqSTDUrHfwBYPiaQWQ7kvOCt9XG1
+eQncN9fZtwRoz6kEw+GGZf1lQ6qtettgobeGk5MJvAaWL50AkTnjgfBe92GDFDD
iMR+FIM91Otlvfc7oXOpcgHLP0UcsTmqGyTXA5H61U4FcXLEzE8qEz7ziZBEKEQ2
+UOmhx11oAC+aQMmZqZUfUan4IELsPn3WDcpOaHnRo+KlARjbtrUbJz1HA6+cqAs
R3rCPGR2kFau+OfylGxkWtj7myqUi5Lcz3+btbFeGseUtPvNVHPcsgw6BNIr0IJl
HDnNYkFK7pCHMqH27auJLpfkbFzC8TGTyufIwf4r/PL00HwMKGZ1H48kG8rz/3Vp
t0Z5OOnv65lwJZ2kgXIYgwd3G0/jCvnJzd1ORFVRfLnQsLhWBO+009EBwbLlqBSU
AC5G8W3J+H43x4yGPQ2tbPXnSc1Aee/F/qt+S35i/Ga1BL3VItje/7/h5OlQa7Wu
8DMCh5NbbOZkBhyKNFjOW2w17XpA+NJIj47RenqGS4wgqYqAab0SHjTpUZ2T/Prp
rGYxRkZiwQpPnCowzJWrmoZdrAIFA+Bcw5y70oWf0htdFNw1OSNlY3QMyGwdrade
F+tyxp9Qjxf1n4v+rkmSDVkgpI3JddTxrFXgbxvSCiLY2Gha0uMUSP21+6dvjFqX
OUqcC3Gozp3LsXIrfBBy1Sl2DsYCn27xkM70PO2YJzvZfQusK3iD97nMa3VnQxzn
aoFiuAoW1JLDt8KhhsmaRACeKSOi2kytBw4TrZWIgu6wbg543RT1EPwtQ/97c8QZ
QgHBl83ZgCNdALFebq4dRiVJSH62b8gKzVbRQmZIy14PN32PHRzv7KBWiw01HSYZ
fSjTiZRRQFy58onhSo58shTvvHDLlcj/qAC5MwNQawSLvr2rJqCqSKZDaKhfY0av
Pd8GSoSKRliu0RKAdE1JnmHMnq0iGyQMM4VqbmrhtAnogoO2lITPnb4Km4KUG7Dn
lhqa55teIkyYUyoPdwEou2PmcUDApR2f70LFaVjhCXZOD6mK4++8UUtgMfNIENR2
zBG5z6SmZMeseANdJsLlorLIChVGXG1VWaZg/8geoPpoVVIwgZg3bldGlklKpism
GCRXSkxkXVS9DPKd5bE6HiVr5pGC7A4yn27HOfq1xr8fFdCeGJyz9RZzdnTmFcIR
F2kecd0BWbwwyIL4NxZI4krZkwFGAUyjAEYMmmbk5mxg4xdE3RE+iHffSdglf6TV
eJzR/X5b1Opa+56hLtJ98+2Hli+7regDcEZqDOmZAmXHDtlYXToJRsxTwbPLtemO
edukfAm4Rjfh0G4umycuYwCDaWYOtGhJR8RXSYX0njQywGNrC2uVcpDVuc8m3Kr3
WHF3vQ9aNXSxc91Cry/iHqdPanjbhRSXpdXhdIgrKgVHOOlQMKzsmnpC6WGLMZTA
AmuWtqdpIfIpilkkeq9OmeybrwgecLodo/XNEonxdJ1J/H0fXS0jdqCicrkO36pu
GYpH5O8UzKkjJOgP4B7sqTaw1ZbwAmwzFmQLNNqUQyOdCCsW8p53ukgTPZ6Y9/B9
x5q5cFO+P5hxAD+XJXbc5oISvz0VKOcabVPOVSMxwTt60az0G4g45Ju/aS/TpTEp
R5H56nqRpMgyG5W4pJ7XzW6DVhvRsv3PFpdEu+JEYDs4hCQdET4NvzHmLWZLs7MU
YahFBLFb/hWVvlgaXNitfMZO/11Hq+eMrtwnKUt9Gr2OnivQ22Bukn0pSpczkhek
iIB8gfwiSgb+QJXB/oV+54D2nf33EpgMX8uZ4rBvRyKyu+LnRQV86QIlYPAHp7uF
kQ6J+m+y6KfKRGf4V6jEVUuYtnWGcGs1/ijUO/Me3R4D3hANs7ZovNCOw+Jb0C7Q
N+OVXvntx6+iQYzULOwop8oDp0n1rXX0x/CbTLiCmcdCgW/BnwE+Xb8ArjVQCLxB
gQK+5OIq2VTvjCULTjLfnXcoeIrerWZFqgOgu/PJ+Z+mq82AnkoAeG/Y1ljgpSYv
E1/Nlf263D5TY88mqpLmZhHDwmVwj56UxwNE/3CXfqLC8nYo1CBN/xe627Yrnx83
m9cxR3xqT51srWMKHqV2vqJyRNWPQriwbnpsSi2zgE+kRmNRY2O2AxEfFBriWTOH
cSecHlu0eAlT61/0j1uXm4LEunVYTykA72FZoQMIMPA4wKdMEOlwXkywJK2LH6pr
UG4gcs2vbK8VYU2LmSwGFW65SvtuWC16yRq2CUhiB8CtAwHzei4KO3kjHBgykX72
+UqsbXMkFBrRRFN4CtphBoDhMT44ISJ3yK/3JNDEPk6ovG37cF9oyQJaA2uHNm4O
Md4gA+3JNrm3rzNy4IytnB+yCl+x+55RD6Lkeba4RbxlJqRVq4Zr/l6ScBAZf8ta
+hk1EPbuoCvHjHrTUYa/qKARmlLF2qLlmSo7QfQ5LJqJ3qUUMTYtoNrXaF4Wb3rD
QEtUJzbE1xXQMIqTCuFupOQFGdZ+l0bZbYtDJkV/IHLF7GMAMyxHHUCwm93j65cC
tLwWFIkuxw5/h0DEHlTFH4ZNp1oRmUXY+wse18/esGglkfYFkMCBEjHARPkHp8fD
nMy/amj1iV8nLih3ZaDGJ5l/jta3YYSNXn8kVnXSDn82l8ahZBuT2OH6w4328K4Q
EYXlUsQHDOp0/oZ8mlPuSie37cD4MVrMY8LUwU2EVcp/x3I3sB6VCYZFLEMvRlw4
VKz3I8JPpgkAJvYoW0107Tmd0k/2iAVkgxRwKvBh0otW3mRcnv/H6NI8MkcoJt0H
ertmc9zG0dJPVOLMis2Q/VltA64TQMx5RYYq3Bei5M9gTx+wPtetO+pxU+uPJFkA
grmDRJ97qEqQ79z2Wz5syLV5l4WsxposPGgnjbl618UOVw3n3xeTC2jeEHnWRaHi
c/zIhF65sjwHrR1MJ6PpUzopedn582fvg/Ggom6I8CbcojWYOkPEtGuPyYhztAA7
oLyvHd/8vEYRoqPF+OqIOROCuTTGaQxodJP9UbSD7GIiKOYgFq8xKm+pXz2k415A
90NKXwPQPN+rURS7NNgZRDgEo36P3efSNBr0qe9zutQzlUWY78Q6J2a0hcz0uAwi
fl6hq1n1n6iK7OW6YXZzlqEH+y9DAbKXvpdzsxQFW3kag+jEMNJ84rOUrVKLB31M
UmWWZdUhNAsnnObxlDKixMuBzoUaeTGu83HdXc2A+s8Qrc6hSI4p5tsAYZmimwpO
5ZWqAptEyS1pGlP3z5XHvBdmpuXWEcmZqtaCv4HpbRa4zFu4oLhbqTf81WNXc0zs
SQOgsH6ISW/1dH/OVJ2EWN/PtBeGOpwVuDJfL2vSYuHveGZVQAPcjsxbTm/zvdIi
Q5J2dlfbuH9EoIsUzzR1ag4lohPdr5KfSeJYIg5D5WEJ2W2FWidgh55nuKrONosl
kUU8SUuF41kwf2h14Fj91RGA7TwAf8PaOaitUe/ioo0Y3s/CQF0NkvIPDiTmqMmt
zyX/HEiH8R7F6DvoC2i2J3pMENoa7eGTVr4+2DjsImwgcl4Tp0x4rRvLc9rMw+jS
/6EvpJe8x6fNAiumVKJyWMN43IwG0uTTwI8/8KRjchmyZFV/jEWZ7joQaXB+ovff
DdVCnnxtt4UC3fqbhTv9mdzWe2Ev49k8RIgg6zj4ysHudQUJy76sf1KOk+GjQh4D
o0xEVStkYkNcCe6Zivhe1wjki4S4ozpEIOEnyh0SUNIY7Tmw+dU7tGaoKI1O20RJ
VyiRB/rvtWNQ6/Jcn+VvxN1qd15Qh1TDmW6l8XpT2UMunfy6PGyi0h+DBkNkjJ1v
XTZIFXNko3yTPRzwW5eFcqth/fWNU4LZpaQosjTofsRNctS76Nn0bjGm6RptLNHT
fF/CTn1xLBf3iv4NMWwlt4YKvAQXqouesCEqld6K79d5m++AEXkYGrFuSs0Y4xuD
BSZveknLwLLTF4zfYuYI9E/slsn4bpzCfuPOm9CXqwDGnrDJ70M9iQW5sCkefhZd
Y0EJ1CDzw3xNDsEGQkOlgE8fKI60vG39ipqQOTzgwplyYcPVCYppfnMhaUcL7LNS
4XiARYr50SZ/AGoHN0vOcoK1R0sX2dh9wlmkutwXopiML6nk/6Vmi4QUTorVDWvQ
NxJ2GSZX+GAzLMf+ulv8n2YqX6sKhxZ/CwYGPIMcZh73vVsWVDR6RShHwfY6VEDa
/1qeOmTD8oV/mTy7t9aWQBh4glwUUFXAq/Q+aXJwPuuLlU+VwrPow2sU8+B1U330
EzRB1QAYXgYjYGPN9HYgotqH37SI66O0nmJ4JlP1AT3VqvLgdULrf6zbzAvejScY
zKwhF0GL8YpZHeZHpcX6IArYuPgX/ehA3gp4AcDnD70pNpkHY8ww4sj/wLDINX8n
yUKlrvEgOZsd9eI/BeEvDq1xsOsufo1yPIHqPmH7ggTbevXlcYyNqmbgMRToW67F
mW3vWx979dL9CmJX2PPO7mBJPfZfCxX1MUyQCH0XWo7qhoRWidggQpoAE2wZvy5/
uk03ciLFPM4twxlrFZ6y1/3Dcub2BMJyO+VDaeBcS/o9J8tV7ppuzOMSxsHmySf5
ka3pxYS6xXmJiZ/ksnSq3ur9kf42mTlXfbPszuxJn8XTlkZXmurdpJn1MD5rph0/
XFFIurMb6dfXk/8OKlshsW7IoPOAMhDB6aN2JUlhJI0EDOkNpa9Qgqn5b3uLE2Lw
b8oKomIFurmntWz1rwZOkO+fn3lCXfXZVWhPDT9JgRf6U8g4z9Xu9LSzAljITcc7
VP7349cvDEv7danwz+zflNhimBRpWRmWdGJN2CZq+T+TcbzeaZfcsuDhYwzCZcmf
hCYBDza/eyEVNw/ktSkxDvORK12jVWqxnsqC/Crl10ME+PJuP1WSQwiQUC61hZCy
iyGO0UT+AgCWn4vVgl/+Gh+xu9kfVkiVxy2XazkGrQsTAw4J/YFP0Q+wGa9jhxBM
svQpdqYTR+PQ3mLfpnr0yDPtUhouXa4JIkbRyAjiDuwhSkk8Ei+Ix7fTKA4RaUsg
zjjCZquX0jFCFwDR+L9j62fBBUfgehfCA9jM0rq+VuxcFKhwk0WKlmZUocsi+uOd
IwoiAJR5L5HlH80MAjMdUgmjFG8XkyBYA+r0E6oPxnwl8pCYshOYp2+8FktPMMDx
w7cp/XeTy0idzUnUCJrauQzWJNUbiHvr4YZ7lO2cIYoBtgkU7gguLF9TxL6p34/8
CQBprFBa9xCUMEF3cWarrY+ym/ekzwmgkQ30Zt7SZeVQ5Aq59SVHJGkSGMmIAu4l
FMTwlVDbRbZkhK5CbUnpKaXn/x3ac+azuJqAKrDIndeHU9slHTpQOeP3EOKw+SrP
pyZokbiIZTs3Ia0Qn1s7N++uBBIoTNEFEmU5QYDckPjHUsHmt0972Tna/ZkuwPKS
NswbUZI6TNCCqhTTy16fEFx6k4iSzsgVLrjyAMdpSNkbv+d3nn08jWthkWwNaDKK
8Ak1hCggXwihWCSUz9Qbr5RnO9CO78Tz1sHmKwJIr2zjJoMzGwZjtAsm4Co2toRE
ezqkBFpWfb0vNFFELCcdywKFTM2toKY3AQ5nRAfHSf3jwMNyjGWnkNRBeNgT7Uxx
+noDsyFzkhv1vKqYlPDls30RckeiJkbJLg+YbyF9WrpyXZ4rRVts7xJawKL7Zn6T
ccyy+EVES/27B+jaU5ISSVc5AlMW2X6A/cCPfLAf9Yv7yDPWEqKQfVAGT0FpQbBW
3Lto4t0WyoEK4SbIW5YfcmaHrG9inBkemDCjUdR64nCsZdtGx6xJsoUEWknDHHoG
NSiaYf26r6waxsJeWxqFqjhN9tnuar1swUv/dijEvZ2PX1ZAy2kIG5ItZFRjDeir
H3yOq8PkxYhV+UjN6nS9DWzq1sBCqK66citw1+vL9/KzW3Gppfz79ii8L9DpQetj
92K5MEiDUmTSyWXcOiHXj1c/6XrnLwiuTDxlvEoHLaKIVUId9Yuh9GCzKor0Vfkq
ePvZY2MEjTQ5tx+rMWWdtQPfrc+yEveuL+WuZPWuCs2TmTClCpDo3lBRTA9oU0gw
MGjV80tbPR7pf5npjJzYlnIg/CtPp7RymSCg0MzIGS9YeuNN7ouNHvKTWoKiFPoW
x+j4wMCtGLD1LNirohMt0m2qS7FNBzadtLcUhZ7uEUwmp+Xs49MTohsiOk43v40J
zvl7hR0saWyVm5fhLxEau/t3kM2rpJHJXPhrKllb8e0Bnu4kP3ZPLTpRwDSZGMOR
DXGs+KqlLGhTK5FKwu8EHgHZNEfLx87DqvVFC3a2KS/7NYMqY2d6XJNOVMW2eZF6
iTokfXScdpu/QC9YQonZ4wmEzxxe6OFbUdU7zqwq6v1C3YV8G5hSx4KxvKoIb+A7
bbMs7ydBpzlyYalMiGIkTI3qQz9x9y1kcslXMdsj1vxq5bihyf/O92rWWwp6udIe
Cr786pioH8ukH5kdpkQBOff7yfAi1RM8r4oAbIRu30iFZdDeEeXpz6fBreQZkug1
JzdxE02WIvD3uQJ2PFqmB9fx1PdCA51RPanAzY7j9PPpA4vCk/NKsMeOchH0pzgv
HsJjRZdIN6XbFbQOubOyhkA3TsY5dDI63AHa7TzJhsQEdga65SR8l/sfbBi+cuJV
f0skA2OqtM1sMA5l1iTwVN1YaWNYtd/O+2pwHG7dfAew6Rizvv6uYZbtrYKe5Grt
9Khg4goR0W1u/Fm68tFUUQTPenZfpaVJIgW51WDtp0TYzKvncI+uUJ0AkjQPqF5W
oaD2LHuxbk9rguY7uTTNQ4/e/LttX7sl3zFkCBuiGCp4aj4atDiv47rN1IaQmL39
vSoIfrLQC2D0vvh+tm8i+LTUvN1F0+IW6lHtPG8k7XRuyDzaOD1IkZCiEAJX1ErG
garpn/oGqzvmAzfu0cydhFZTb/ZdkauyxnEPyoHk0LzDQWtuhJ4WVHVGQcK4lKFj
wMltg8Sy1klp05N+9hcITfdxpQ22NtbPsLMU2ASiraVJxoIEn6e30GkjfKEW+aGJ
dROVZoodADpIPiUjcqVto208fKSITsDXyJnwZIUCHLXJ1vNbB7Vv77G9LFU/2n01
SFZeZt1MDIskwoxT/xUI4gGZEPzg7RVZH8Ur4G0IrBU04i9UrCSd0IBhh6UmO2fT
BnSTTUvx8YK+x3L5AjHQPIryi++hauz87KRMF78x6y+IOAnTFW+cpGk35mRi1ON4
Ydst1Z2OC2BRjM2xbt0J0v55yJ0NznlFPSiSzD2wuVMaiDyncYHmnCkIebJcW9kz
QEN3UNcUbxkPoC2wnHsPBDUEq5gis1brHwqZNrwrxdphngZpaqn/ImEk2dAVvJ1d
Vs6CSkE/uZ0ZtCnoUtj3ltu8yZE5Xdr8NPRVy4T3DiaQ0Ml9OeAnDUeKUeK5xpzw
ZVy4X0SMcDM3SmBZPYbfOkDYNLabT1m8TgbONIXan1Jz0GcXopAotOCjHle4DO4s
4Y+Fv3usx3Evm+T/JJ1zXkQjhupoD/n8aX0sOW+L3e3rY8sa2Pov+JozeE1+5FR1
DC7dQyak8muxbbd13k3ak2DIXua2V/doAvuhXFGou6KTkEqPpIXWZRgRt5X2Zlfq
8jFhmX4hxYv7lWctDmevcx9bM67VmYYUKp33Eqiik7AXMrZJThgXYnR88SGmd9i6
XmjvZWJfPed1iXOSurJq0qiQh7YD1q4Z8ho3/yNhobDIuGtGUva0xwXT14xsSLvQ
RaIRmW5DvmQixx1sQn2NcEqdipoaZlxW5BR+HZ8RgQHslyX16UPA4wnzKzAI1iUR
w0fI+Dx4zeBxKZIfJ2/LjOjHoVJht/uM+CzLxMUpuFA9TceInS8IkE3ukChzGJTb
fiGOw5HwyHNiovvj7IbAKPqAxkP3KSkkQHGjsDFpwPgWsKKgVWS3bqqczpRC7Pww
bC3p1Ewx2OkkHaapRKq/EUvLbdyq5Y5lKqGczVtGChNqSVVK95f06btjvoqmbHJ+
SBkvtRKzkE2o0BkzUsxdXpXg+TNgxaABJDlftZKeEtNSW69lbYj01xdNWu70h+xP
T6TfnmMOxHXmamJWWZmVVaExomGUyNh/WdP3hMSrNYecK2niaG3NZwq+rYBAiYjM
rwapV0Hh7acIeyom72xr7dz0Zm7NUllbTl8UvY9+ENkkzy2y1tvYpJOxZgwJcKwF
I5lreljLpSNH2/eZ3f5fKi5KdVm6tnyCsCy0ns62yhPr8hnGsuU41w2kjaJy0erk
9tAMSX3qd6EyrBflENmK+txsRZRBoQGdpASZzw2uHu+T016Y2PIeSaJtm9IAknzi
1YK7sCUzvpdzGWGPJtlftsxOPkueHxj47afvT9pMmpqNo4wl5ogJPDHZvv2XQ/qF
WLq4cxYPh7Sz7F1SG6S5ibIO1DzS2McNmWVzf8zxJJ/NVmHzSPKNC/iXp47h/5qM
aUZkxr6KBJrcKUyrutYZ6GbGjYUrXTcJvTZ+EHPI5Xrwga6aNexs1rUR8w5gwYod
DuxHh1nhwuXsIh3RckRQzpZDZ/mgNOsZZCBNapCxs4zjVSGSbKxe7gT/y8fPhAt/
CGak/q3VBqyT5LCDXoz6hmslV4wSDCQR3Itw8RdzfwNxXG4RULN3by7XoLTubEsd
ZkEe3MH3qERtlO3MC10zsgDSC8efdNiMhpGQTVpUZUbw4/ApYA6Z8jvITZIHW3ma
LzUeIlGhPr3Q2veuc1tSR8OzUjyilxZx6oZx4LKs/3pdKMSXUbcdJ2hR8YQEiwuI
nQ9JfJRj8czGgROKi+ocU0G2aFPufeXqly4b5cpNI8UInrk9kpEBpR/1IgM4IfQY
4bSxLBNNyV56gphI6phRZtIoeZHB++IgCqpkGOl7ShqepGBuCuoMk4UtzH3ZASdw
xrkV1+Sceu+Gl0NYV0taYnLfgt/YOzaLEcCNetWr7EZRTqnTPNaFVUN7Ct8BjH47
evm/CDd9bg22ee2eaW2mmblK1p+96/vBh8MtyY4zxO7C6DOXr2RU2XVd3QHCGmFr
aXGjqUfGUFQR8sGP28ptA/60eO6Fc+/ThZlqPSqjgl7n7z/MFmh5ElCdfIzLkSlN
c9i44iXjZQxcWyT5LTAVEBA6JS1td2wYFa25LZ5+VZHRCxX8V4bD7Gx9OeY7+g3R
+7rROeZc+N/u4mfe5IHZbcooXffC5toO7ooXs9MaZNXzAOQ7vl28MMyCJ8/GEHQ9
X0fSTXKrH0TaYWE8mPID6xo7H6J2rvReNmm65fCj+Cd9yBM3LkP3RSz+mHqXyN5f
1gQ8J2wc9w8rdc+jAtPCOYi9Mwc7Y2ATJRrK1EbtvdO3cDghEAAtmtMnYIDiNsxi
aVutDX2GrVNyvgYoWVP/VIpYzSk68SbhOisZyArwCNHZTANgzOcxHdkFFNX6PzOj
sEIDKmImaeRBZA+EyUh87GPLvBnI+J1OXUSrNpNxWaJSA+DXmsPMivWL5HMmhjsV
61S6lQE+S1vG1rCNlUrbmYM9oyvS90D7ZCTY5rxYds1IRJfnYC0MgyGje7HFFTdo
jHzNrh6csiIJV7x+k5nXfXCQsmXnoRd8Dnu4XIvwTCYwiACQHS5MXDNlgX/H63zI
gT/diqjsFeiZy5OF/zT7gdHDAR6VW4Jb8Fl+93DTvej7Rb+E7Qv6PuiRRxBMFAMN
6l7+RCT0yU9hLsjWlpvQpjbbOuaYYynFJ/afq8tbsZKrYLZjIBgtyrFQqNDXc6Cl
eMoJoxqTBvwvUhP2ZRZgLC0WTqOaWb6TXLn9W//opILfaPPKfV3gXtj6SX6FpDs4
SU2/pLEWJVw6yjMjZ0ZTP1ZVNboUXuT5zHYU/BU2DNOsT+mCPN+39BOytlXred6l
aFmFiEpnAl9eZsA74i+aDzRakljE+t88QhmhYII4vow8PsRJyNevSqeXfW1ICr68
kkLlhjxlqOqHSnRPFKIQ1ait24fb0wOaohVw9MSRyzWYZkqN8MFrzrUDXxdgnmgZ
kg0ItTuoMF3FJ5rt/qOEYyGFdBAuaFDh39LgLXLASWA3BJmYsQP85Hl0Gjowt2iw
wlz3nFGKEle2jQLwlFG1JgipV2c9vtpM64q2QRvZ9zN9lFF8YGtRIp3Szs+E2w0l
FvKRkjpCDhDCf78ad6mnt10TNote5u6GahDBUuM5B0fQEWwTicqdVrhZOUAdbqjf
YbG5ovNeh2YfFoCFT12+uWXyX0LpXTvJlrBrzYuCyzQ8Rh1hg191yhBn2nJVnKsg
ciuV2d3wjRwdo9Knn3EPZU7jP9IwFoZic2pn1f6pPS4IbMVB+a4quULdDs3pVMqb
rzr8i2xUP7Tcl9zdjducdZIRFubF5duRILf6Tmyh/zOUn6TK8fvHR6xj1nK0T6dL
Asnbv+fYfDsA5RJed47PjZ4cWYqIO26drkBPxR8EdGCF5P/FsBCU/2uym9rssolr
KuMbUju5VsosexAE2l0HQBe1uEY+xzjcmEPmc6IHxb+igjS2v9lkZ1/J/UyitEsG
qQzxXde0kR8nKQFuLk9KaO+/smytCl9fLSBQPZfY6IqID1OkpeAvoKeXcwBf8+zA
VsJAOon/S6QugLntMJRFFVyj8ALtL0uZn0x3zZ/xtn3BW/fdthhmC7AisOfRH9Em
G0ZQ1LNb6UpjrvonAG8cSJlHLui4+ripAvckfB/6CtBHi1GuqSwuofdiRQgMnl10
K3XpiBqSjnfNUDX4BE1LJMMf6GMg3JasAtTgo6dI8EfBRNlGsjPHcTldbRutw95W
CgIq2PYJb1Cn3Orklm4OV84RSaf3pLArw6Dj69X9jrtrxO0BiWJw6TPiRsgX5v1h
wEtbfs4u2oUCWdzgBwmtIWa9DlC/O4R+gf+pPcCffhVnaT3pmvYD808HwMVOnmap
1xuMe3Ozm9f7CSGvTTKcTu9uHwP9619j3+rTDEBg/ROm8c+cqmW0W3e9KfVtFdh3
ilCXkHLNZl5DY3r8gMSGXk/n3IGqFc2Ttm4JI5R7Jh2Ys3wYzzCpm20pXjBXVuwm
MIEgqIu8MFTkfb9//E6LwAknWVl2PK8zpQWQDw842gZJ6XsaYRdPShhd0+n2gODw
nH8+7aQ3YxpR9/qum15DzrdYAxP9XqCJs82jVt6pYee6IYjjUV1bPo5F2aFVyejH
htaZQ5W1BZiLqoQgzFio5mIMYFY5s1TzmZoc7zPkigwVd6y6LwfviOX+C8dMHMlV
WEJ7H/a36147wG7oOI0vdW6mnNSE525jFvkcGpw47y6uGuGamcBKSOSG4jfRuCgY
9M4o0JtqH4hlK28SJGfaEYl5cWIOF6QprBI4V5FbxDDnnDxIEeLSGR9wlttXNV3o
TNTTv+1Ld08ZsI7IyUB2McSn2zYh2ppO5PKTi26sIAutX/xCY/HQ1r4xBlFo6O7D
YhkPKroW/U0fMAHBDoP78H4q76S0RFYqKV9IeIYq0IuPZYdycXoDRV4gkm8azLrl
uf1ouIq4btLOmcz0qx9WNBdR7CFBvXdyw8VA5mc5l3PabXmw8xCZdA3yFp8S7cj6
QHs866oKoCMgGTKdH7qd6oLBI1WIyyUjenQ8srv8JhsIiP7U5N5hbB11A9l0bc9S
ZW9KBJZOuVDOGNtw5EUN1GyVDoAn0VIM/yhybtUPeyT5/CGOC3uH2yC2YI48XlKK
RUaHSeSuhLHGX+ACUUR9uR0BjjpUTrAS75+rO3rZDvJhB7p6pkAiKTVdmr9P16ag
pASYnQ97LQM/J+wPzakjqLokGPEKwLRe29jT5GKy/t/D4vavCAvfJG715x1AA197
guldoWGSvaU4jKtcykd69q6pGTvresHBQ7PkE7HZ18E+rLWipKvUQay3g+aAN0aD
Bk4+n8nG6uWEvyLZ71Vu6L689IXq61akv7XtPuIBcGzR23kalK+NZ1C6TMBrgqR2
vAVoocxeksLqbEzcXa6hCB2Ri1YmrXfAybT8JOaSTXCuIGcChxUHrRNJ3o8pySL9
ENAkRpQQSrAMQQRNTc9ufDmKMmyLqoRj9vlsB51CMMs57A6osQgewfdbBgoDihsj
sT0NZoa/YamvO5TOCbx3DxfhfVNiWv1amFYGhyx+/I+v4pWTh/JnJ11m+z0y698K
6TbM4RepgziR+mxuYsrciuMHn1CBYPt76nq+WDX32/n663BAYB9gFmHoVY1xpQ70
m8TEB/D5cnIo/FOpV3gwI14fkIY4m4nDupuhrah/jJtkc0QtEiMhKgWud/MrSpLT
7GWHsA6S1V9ecVrS6GSMPfCNCjErCjNBjSEKToyibPh7fDQm7q8FuXjZtZl3i/sz
56Qg8M8YBHX4pcRJcNwQ7//RaidM/7rTuX8QOSCC66PP+L2u9kIIxauhYCylF1Xb
KuIUV7pk0eV8vR5pWDoHVg06NTWyEt+IheKiI5UDtdzoBWXWRT0B+cw+57Mp2Y1O
y89YVYNm9tSPQdGlp1IX0iTnJFqGpJtS3MMYK5k7s99n/FAgvT8fhjT7OddVb+Di
tv74IkIzsO434ggcUvFMgPlPlyXMwGRpCpcyR9yeqvJJFoHVuIOd6PhWzt6aA80p
78OcZDvTJlHJQnazHcjp8c4aNTReGgzU/Uk/SrZb9WS4S0EGM6HWubNl7Xg5lJxn
4mWQwHZmEsCA9yNsT9R14QOTrqFUYDmtd0vW9eONCS7vmVG+56LXZu0S3bdCKkbD
LCcRTpGQ1u1LTluTW5CWyM/7CX4eieyYmqhTYM9mQKnzJyRXsq+N/XsMyoIsmNyH
qCJGkzWZd4oDbKfe41WBIvXoMOw7+XUXVOY4fJpP1UN3GjxGWWcQjRUcaI0OPZD8
PkCtqynL8c4m7/UbZVj61ZmJVpYU/e3zY8koY9Ms+BMZC4/IRMGd7WiHxSeqiB0E
maoXm5G5nP0J8DT1v80GSvTlVZpq5uB/RZH+VFyTmH6Wq0aOdxO1xck8c2vQ7OkH
FUC6NsDmMfYyu6uQmK4JGCYJYp3UyhdwjwSLMbXtACBlCXvyiRRwH+M4Aa6T8xe8
ePqOFzvUT+/NosVNYc5gEkaJEEKTRIwYxwYYC+fd8XK8Ep8Bv1xZVK4BrET3gsTV
vbwsdpLSizWmr9t4dsbqAnvGJOPtLvUs6gBo4dhVCoRN9kA5J+xlnuo7qhURqvsB
WY5o7tJbfi7BLkhrstQzc2fVSQn2FbYK7uaOTWwOQr+lJUksxZ2kDL0yUiFUDXxu
7xyP4qVrI3DAjoGoA2dwqDnEjEnptDurf/O+OL8yNsMZoWtWgCXG7iwFBvar+ZZb
cfIPGODlEHfwemvbe9tAufQn/V3RaJARVTA64HOMAdcA4EwL+vF8CqZc8VSL1s41
52NY2GCMm970VZoFxgEv98MHgLM0E5Fx2F5MQn5utD78VMc+YhRGGhq0iN8mmYoC
L5FyIQx48LmxRM9bOGLzvX4eVslT6s6tFGH0iGHHqpzlTBomcmdkF9VjzfOwabBQ
piuC+1SS60OVsHHp2cDizgLjYyqtDh8SovY5kxNuWLw43WWc13Pa8uk+juvlew3p
7GvDR2uKc6npF+Y1Y41Wg0DEQw7Pd/oRvWaYh9Go/oQauj3edP525NjV94NZOSTS
Nr1gxyjQUxgmiN4k5N6I0sBeDKdL5UMbmq2N/zLOaZkT0QpjL9Zhhur05plJbZfs
bdW0tE/z8mnSgZron4/AKq4eyS+Z8jCd8oVWq/iCAX/qI+41iqY6pkYL0N8juruM
4jUF6bfEsrY0GVoqAjDSrj1TTM9EN41vmBbaAMdg5Oq/stmi1dwSIwlAGLc5oa5v
EP/fGb7PwSldcglHGFvKlWFU+BGhtOaOj5BluiMPRPN+R2RqM/6MhrOVAM+0M0JC
yuQ+w3VOg0KrA8EZ5iMVJ/sFBpNejTZjVDT5XyBbkYNDNMD3xxqZc+jqnkQNTalV
TbtCmi33oHxQe5FrWQokpwCfoF/pfVBZl0ksO4w2zC6yG6/RMu5rnVi5Fuhv46jG
8Y0FqHl+Sb6HR0D47wwX24Ww9o1KsR23i5GNiWc+C4ad4Vai8n2zHiRkTRyIaTCv
S6ktySKtj2gKZA60w8ksofJwfI2YWRnpNdVv5nUI8j4yWi1NbfwmLBreKBJW+RTQ
MpVMcvLnERZpu4jekkiyMSjoTxDEyjNDjuJmmQGMMuqeyWD+GsZVIwOhSRVTG3Cd
Rr+UMgEnmo3fk/xVNGcYuqwlLFU69UbZG6r7ZTkfPJcMesGMvlmRmizIuZzBRlg0
B4v/qz5RGUfN3npJ1mbBLLaJHxojXzIkFQra/blCghAGslw62RLpeIiktRqN8+c/
4GiJV4XuHxv/eUaU03yDmFLe1lm8k/5ZVR7NQHlN/BBT+s3X1Oy8+ilLS1jvTe5N
zcEWHbVM93+2qiBTgQiLRpX6lGopGk0jKM2VM2jDkbLFgsSwT+LP6Heo01E1IcHy
CIyefzYLLiWWY5E3hrWCZYQbZjH10mf4eBwDmRrQF3xvGTbGtKd8sexTMGzOb76C
7R5XJW3x0boMAS9O8bv57ZD/iaT9aQQaAvdjSeFw528VTDeIzE15Y0BUD9TrhKMD
0XTFpo0+LgN3JY1lYMqJ/lOVUikmYx3T53JcA1NbI0TVXnISfG7s3iUbrrJ3qQ7w
xqMTEk2qkQOMEaGwbAIL+4GLTNYSA4//yigfwLYLW7ABsj2/v+GaS58La2RNKkTh
69n6IV+bWF20SkjD68ODdMTixlMkNPGK8ZEaF6MTVOrb/9PnPGa6QCvBG2m0s9f2
uFEI3IMS+1cr4aDnavZo0SGIEzRs9ne1ULBt+eC+me/3TK5/m/oeGsliEdWWkiwr
xlQq4gAyOS66AOMWlLF/I337Rb7rlgPa8OeTU9A1IcFL2oZ2tPxm0CJ9zJJQpbNi
hxFUDVAz3pwDjIL3OZeEvI/3BKhkRcKGctHBhwG1eaPmYzFItVYGkOTdTHTWmW4Q
1oJxOZq8jh5s6f2ZTIexxGuzujXzLhfrELLkSRHg9csKC7XZo4qzjPD6/566bquY
ebciyWh2S6feD8u8Ph4SzIkYVHSi7Bt0u+1YXIHOBlxslRUOdjDywZaFL7qapD5d
7Vkl3+AnGWfoeJcU3MRObXT5qRDvfyxvuQ7G5D2NeHsybmnOSHXdltOiw25mpzC9
XRqHv//xxjfO/O28Jg4EZ9NIno7pUBZwTbXz447NRCTySqwlqxOzL6qXfyXlyuhD
apyR2NDlwxRVA7tg5fRF/MlXxCx0/RX56luF1GuoMii2NHajEg0/I526Iq9yiA48
7Y6IiRfkRRR0ZdWkunp7Dzcy+zPFacMuUrCZeU10fMo9zfq8N9nzEai9WM5cMeTS
9VTZRraGaqKM9TDLJLCjP59rKdvEwfBL62gFgNJNtSgwJ8fdZA5OnXSTLCcjX9tR
vsGYYeLLGTJMB39w4yOAN63zxGNEzUmmOMGRd0a4+pUzjcU+a2+ONlsfcHMosXRQ
5AlT4NEyrZAyYHrVZA3uKO2YdQRpHrWIhugRRpLjF62NE+bxwLoaRNobPyK5Sa6l
WUpNTlvBQbVBqNNE+tbgpk1lKPDIelADw2SFpwK2IXElNhmDh8q+jl24m1M/PAfn
ZernS0+2H/OHkJFgcw3KnbwWzLQf+p+kA7NH0VGsZgsMAa1uhj/mhXOm8uOWM18i
b74JljtIv5ZMGVNqVzigPK9Pr2PiNnqWUNpxE91W9vmT/WGyMC30TdAiv6iN7eYC
h67j6UnE4CmCXrtvjw2YVtJLux7fqwv4n99eQivlBFqLdRqbdlOJJBP2HtPlvEkF
BxnmbBO7+kBRsJuM1bgyUw890FqgQus7LPZhW5F4SwT6XOKz3dJ4gzEHPPAZZlgI
adCbaq5b0tNISBjdGyaTaOCHIXODFTsdF1t/hf0SvCj7s2lGCVXDQitxyGwazDON
tY06cS35KobE+NpVHFL1OjNQ58snXDo8inS07uJ+5YM3zOm1kWIIACNNc3RaCgXR
hn54KtFwEmXsVrqCbifJMSGwcOdeaz/SBHkdxXZJE4DjXMNyMMR37UbKdOg0p5I+
6s7K90+2ilKKdb73JUED8YUxl38PpVa2LFmgpHR6iX3E/Yt2jzWATtdkZcpdf3RF
Yij7UqeaZEcNf5PrLLLiAM7BbVjCZgTQcQQDdZcq5Jj9/4SaLD8NRLe1CeuE3OBf
vb7/jwk4/1CPJe+9Zd7ctTfum8OA6IBSv9BemgHJ3tkkhH1bRQr4V2CEpDoAeuH8
DOm7E18JMVLKI4GlDZXMhtjSHV8e8bHvbM2JaTfM6J/WU513/qEZej/eXNE70Am6
XXtfbyv5NS+3zqNj5MgxmiNSa4J29KaARP8cC9uOFyWHRjQxt797gSKmBRcCYPwe
V1zfxjfewAUW8FwQ2Unuk1Krz4XjsPvPPZ4kv/MJNCgjE4QKIbqivNFZSqxukj2k
CG+XZhhqPktdAmaXIb+jbM5T28yJoYTeImepGYEiCk5KRY3NK5uRFNeNn8Wuc8qB
TTsqhfRJbAxpcLJV3Hix5bgTpFc5kCAgMYC1tffLcwgDU0Oelrhtue0D/XYd+MVO
oHx9W3e+MydbEATtZG6njj+TfuXwTSPwJAY6jSF54xFVWI2/G5CSpqGpG+Lw9w+Y
gpNzW6lyc0S0vUgQgnGbrNfQsKFTx0UT85uMSPctfWmRMVOS1HVQ+Oal0O8V6MkZ
XRL/rxQNkF95cuULa/m+QSk3OrpfreWyC6az9q3Jqbcr7XtXy0X0xIvQZHHl1Fbi
N8VTqdslz5txxk7TDJCVLsNz1g96fRCtQtOK46jm/p5lUDFucxjmuyDPQr7py/Rh
pyBAJ9o941anje5/bNu7u9xyDDRn2onqz73l3RcjdHP/JeCB7Kx7lIC08lh59C1n
S/StbdJMZm2b7icLS3fkZ9xthljRbqCxetoWj3F0Ab2TxT26kjm/+I+BeH8X+uTx
iDMImNjN5IcFy0mcNy/06Fk9NU/Rou/c0oUHczdm4HKTbv6xqvJOep+T8ml+8nWx
enQ1dRvBRutmbVJOcKIgoQ0vDrE1HFwzkt9Fi25ACryZRU3U5nFelWNUlOVBuZNe
9bqOcbFWV0UTbJyZdvMFpeHXpqv+5nFhySJsY2PnmqjCwgae3R3x6e0INNPSigPl
tfEajBYAtc+XuPtSwof0A1ENdrZxj/ThxaVfX3sP69SmhaPA8BH6BKDMRkZiy5mI
rrUlf9wXEfJAc75NtA9sHvQaOdz6WULLvMZKs8tipsMyKtg9l87r9OfAT2a9ze3A
nY7MHpQBK+l1XBnEXHFVcXFSt+6/YJUMvSnPJFBJIuaruAZlQwSJx6845Szp0NRz
5XuogcJY4fM74OHfmTB0wSZjZx1x5+3As2lMhZV8nTr4Va2c7Y0yLBkB0vs1kbhD
TvKG2M7fPS2MBh88hac+UaoNxWJnQIZmhX6Jv39w07WY7Dji3B+D3SaHzHVxfbL/
v71QGPXG0U/ubaUJidn6c6nEP+oSIyVTAvnxXYLsdaFl78EZZFqmLB5cdyfdcAMZ
OWcdjyfnIcYvyMbCOM2z+w67lu42DjwZ2hlvtRN7TZ6qIAQGw7kNqW/o7o5rgOnO
9lwq0gAjBdo4V357Tej3VyM/Hty/BTXDGgwD75lAnj7RlO4u9pAKOafZQ1AuOAzr
AWfEK+5IcG54HvIx/qYqQknp2M07Q4sbVVlCSOKEyFITJNi0Axz87lVWyctQuhXR
DXKmioGsQLmA8mZE0hr2SAhoYhjYRp5a5azTh6eltwlSybWkNBx5NQRyphoLdl+a
b8Q2EGM7hChR1G8+OQepPKd13tamS7c+o/QW9M7Iy9OD7QU64fvf/cs1SeAP3CVA
Elt35GyhJ3GVcMw72mlDhMftF5ubhlzX9qaxM9pjqUdbADVUXpD7JwqvJkCH15Ks
zv+wQnnmAZ6Qr2T4amL8zxsD7CjPYe4UKw+BjMEVZ8rlmfuWkRszxrnieeog7TYy
ELv8GmWe15wDiiawEkqJeNXj73m79UT6eAXTrSMlbBOGyzWeTHqkVrB2DJuBZp2f
uuI1gdJqJQPAfdWuCpeP3hs4v3D2Sm8G898S67sTclQ2Eke1MjCOmH8IMlT9yUWk
gi3NnYGMFy7w1xoT/h+yqnYy4UqRi4w8pFIaJUrp7/uRE0b9rHBp5Z8VvU2IshTG
1T3kEqyD95e0TiPrNHc28TrL+r+e4bCSnUeLAuP6o04NIbEO50W768rCjU0wnBe6
ZDLXI/Y/WCy7DxU0q6AuKx+ivNUuibxXHjiv1WSIsNkda6O6XP28tySBjtF7JYFE
sqDXOc2JUBZYYKNhiDwoXblDql+cBe8d6zQIU8GLASnIv2hM8INg1xOIhCyWK75s
I88eBCW//UsqytGC/Fn/JpOTEs0gsDYDXzLGqKRqbY2eqd0Yn13+oufVr7FUErSI
KHDPWg8fz9hl3BsYrmkGhNNsblh0tyt1ZpikwvD56rtKlBzpxFOce8m5VYCAzx8H
l+6OZFGQo/tz/M80G3J1iQnOXfof22z4tqLa5ZpdD7uShe153si3/ZQ0Yvu6Sv2W
4oHwheDQWXB5C3ommZe8a/DbfmkOdafQ4KIBuDfVXocEVF5aF0X45C8OYRnuYz2t
ZOHTdgm4jnoIzE5ZuT6EbRbATjolgDuSJ95pYx3I0MizAL62BEMqDSQEiYzzCclR
LFX+IqVRpRptVCbtT/TXjQoeoTtDx0y/W7L2b+RE4AlwCSpdjMNvsWbHEa/gc8Kb
MfFIns6V52MQGomNjtE6JdzS1DGblueddVW/YgsIU9QfKe5wfnhHidqmuBKUWkof
d2rnHbn3xSlIo8x4ru4t+rbwNWe1YYWY2iZsLGMsCAAQxPk5Jd8YJeALaajD6F0U
4po70LaJD03y0x3bKCfdO4yT8YQ7wrX4vRfO7QIqsbMQDqHGQBudP4WpKYCHKLP4
VboBk7lG4uVJIK5uWuHitY7hVWs38BaW0sAi5EC3MMRnfifdgY9dCRI8wD7xxa/O
Gl3N3hQ98bHSL3qRoh/bEBjGpN4MZZgb01M/Ld6sAazWEUPFXb8aVYGnCgww3s6r
Z8QKXowz+vXLhLWMyB9lRN5lyqZz3jCErQrDeZSZj4y/86c13hv15QTIJHLu3kYc
z7zae83v25TtniZTNn2OHp/Hq3IZ4xQh4u8zn2d52EdOU3MbV/RRRe5Oe59fjFGv
qcMCgzEc+uBEn2ff0dGCBbR8ORRhDUTE+4lZoVwwHVDmnleOfjV0j+SimWtLSk3/
99kdb35bEQiGzPHwBLNXHwpo3R8jY5dl7gdtxBNNAwovCWC6VeyootUD0ujbQ0rP
oxoQ8F3F50VvBuezoZtTPNJu9WPufYrQ+5akXrSZQbQGFe4uzP9vkAllMxetrJ5p
kSp7tFowMxMfpOdgYsjLyf2DdKKKRwi5qG8OsRjj71slYTq7541yVU/1eMCKxiNa
epOAtm3p9jgkHZ7yWhmKwcS7sCpxRlEBdR3LifO//1bnCqUGJcQ9YmJ8S+RBQVly
4c9hbXIA2p+V7ekVtD6ejbwu37nM2uSxm82I2GS7+BWk7ted70mGxuOZfSfLD/8J
bN07+mBiNDdFkOIwFl7gufGnM75TmVWl6YtMnsNHaSFRBdhfSElrvLtjysswYfQy
TX9FvCwW5O73qIwTnzl7CPexJoAdRIIPPdBx2KZzMF3uAYe517AcKj8PZuPPNLkz
QioTZkfyiWr4kAIpBRT2dj56Y9e7IXxCGFrfT30ucuSkBE6Q7c4cqtA6c7YhIKFF
5SZcZK6Vo23ayTVd3m8uUxljBYkwTKxPdqppGyNjfKs1Dg/CRDpF68vf0FT5O6P9
J64ReRFwCInZMlOslTw9bAggx+ni1pfNEpS1FiPynU7vyUcbGENLw8dHfWT87Qoy
HyouooUpQpf4HNuLIm2thZMoVEiOv1rDib/JXUF6Fax6X4mfaY3xQJOP4+Pf85Gw
z4IpuTiSm/aVjrChqZRUhhl8FiCZpggsk9K24xSz2vL4lrNBcJED6YdaZwCJZ+BY
Fm/MoDPNZes7SfJh7Jo3+lsls41ru5SgyG4nR2UUboBx9ZaTXoLnt0tUrTCQr1Vj
8wYm1m+WvwlWu2JZ4fWPjN/TvUiffbFpaeDyM8DpkxQunpLu17NoUsucNLwM3d2B
zWSUmOlAQvUjh37eYuLMB0ZXoyXL/hpvb4XPFFSNq7frENyvSP1oEHFmU3o4B98B
/k1/03fJloIkQuw4ccQ7Y2vb5Y8MQotKz0ACCNWORRKMP2EEGM5MYh/LxFNDZoaF
42ne77lh7wovmdIVQhYeLsMnKB3/HAmLPLx+1B7D3GjPCvmHVD7zRFJxfbaE100s
7ZAVAI8ZIQcl+e0pW7H4KK0g4hC/zQ0L30lyi9WCp3H++C6sATBenNg42YxTHOsc
5O3z5HIPCQVe8k0swo9EqWhzZGkjCZNc5isFN79V8Ow5SX72ivGqZ88NLGza5W2K
GWBF1ITNJ2yMG8x5dewKWLblx9K+o7obGNFS/h5qVtJkZd2HsLH5k6HeGXZSARZ8
t3Ir5IGH3aNFrKlxmL4DPyFcoRBMdHN+v4/7N9LlscPkaZ46LUyISh72H6JE/Tqm
uB05Yt4vusxMeI0PTp8ZILEkVME78YkpCfwt+/4dNjG03LOIYdn2OUn91yVt1R46
7Vk2Z2ROAE+Vne2UzpdmJoPA9gbXU53ukBbOnST1+QEuNCU+8PouBRxilMmOrJjy
xaPnR9/lKgJmw/tpc9xLJ052+i5QqJKDBhO9LIl/GY5tubwzGVAOZszRt/mZnR7s
qyEOTJAx5fPnzKTNJcmeikH696ratNGcYRzEPL3vC7toaC9QP1BxOOonqwe7gDNM
tHClqB4JVxLGfDvUAWBcYnto9/KcuV6xqBThayO+MVlL8OckRArWGJ7JSE0Adr3N
2bvMoHmQNfqBeTw3r6rfDkw2bWdaMdMHY719BSiJ8E2UOEehunqrgNxszdjOonNU
PcgsX+zfBupsworqNoq6YPFQWk6KS7BvPquubMengrEipsGtUcPb1ywaM6+KUffD
kbxbP0KLvDuRj2mUIdNgbz3pMf4iqIkVZ5THyi7ZkVqH0KzbUbCN8EQTJETxeTVH
PqJw3C3MOOaszMTb8xZ8odUv3tU7AsWmMeaz0atZ/zb63CmSvYyK85F2HQXC28+1
8+/0vhYdWOgU+NyXZTd70MyWdOry+DGzCLpn2hdANVUQKmTBycdjFQSWJN3gDGui
2YVs5r1vveuOGLcyMoGylyH5Qfz4EbLJqu6MWGy2Ek8EV5RFiiW0wPJa52e+AfKo
233lJ+tMkiNLTOxYzlGZm4yAO1Kvfx2ADaUbHX9BPt/KV1MwS0UtfMFL/+PKIUm6
RmTgMGR2b9QDf2aXaRkCPMYqs/X0ZKjqGoOHw3HrV2Kulr6klZOPJleMi1GPvxOE
zYWZox4MiqTA4zkS4yT1I3uatzj23os9l6sa9abgordW/SY26CL6rWCMsTTAOp/K
f5BpHzNGn2Jf930lUORWCjgSv+oHxUEFef6JMQYy6G7xnR6uCD6PaWzpT3JhObWG
eCGDAneqj+u2hhemiNFRAsAOCfgzwh0lnMqllQiHVr5Fu81I0A3Q66SufV1VOrf+
GgtEclGH9OT4hIfywC9zmONZY5zGxiczSOJrtP85x6PXRcNXNUabGn9gry46tizX
B64iDrmxgzD4rQ3n10mCZpGTuKM/Uaw2TQYXL0A5kQ1uTdz7tQ7bJGkktEBnTy8U
JPFWlUZri8ch1MJCrLAN4shZ1Y0OX4fk+A3wgI5mDpme6ffK2SY+BGJ9+uvWIKnJ
0kj9/e2c1zNWFXu9vXUKw7I38zZNGRJ/QKYZtrOlzAURSeXU0kJIKIuZUTROcuqo
wLVplv7iqIjGx2+pJg94jmaLYZVYZ/PjLGXzGyp5l6IchgFSw6/FzMy4Ld0jdBvr
FnSJw/jX5kVtmi73vqU/VevBFO9JM8Ll638SYCncv30RC6tJeJ8+GRCg1DT7+x5Z
5NVVGZ7jQVXt59N70qGaPOH7WzP/hTMrjCvX/5EGWVSfnmUQCOMWS1SZUjNf68ej
R1fekh+f9r6m7XGze4Kkzll34C34wrxSvdGqaXcWm+LWs2kU9PfnveHnHsVB7xuB
8ai420vI1iehTvoLq5gDCYbiR1LlQCSXVFGRJfWdeaYhAwouWZLDELV/XAWP4CNS
nH2+sLlFC9HQ76pwXKAyfUg6P6kNhRybtc3TpSAUo/tVOSJB9VoHLNI/mFPo3vjZ
S4BYgn+8u2nicPmBW9j5rgArnufuctsAXdP0148rjyCO7o5gItPLy9vXuSoV/Dgc
Z8uRfoqAYpzSzA9hncH5IYJ+hXPBLeVxdhUfKV/jcj9m43kbX+DGllWiF3wxhMYr
4ppMdxsuIakxVs2Jdw10n9QIoTC+9N2BrKv9s4ak8Ir8zHrNvEGIncue6S4FpTW1
zLxqRwhRZva64egqrg3pXobO73itbJ/271jE1OvepYjq9w10n8Zbb6VGSykBLcFs
UrFaV3usgELZPOI3QumS9MyLyqDqxiMbzfuuchT6a6L5Rwq76RZhtmnYLlcp6p2i
BCdT/nAIntbTCnOGafq4DkBPfPUk+eXO4JHMZlphR8sTPCFowAFlItI7SQK7NVJv
bQIYT6xnbrDKIKo6zd6dlmQUr0z8IxHeq4nNaCY1uYluDw4MX1Q1XWeRBVQvtKZ/
Td+SQxpbJ999S6UwU72JorbUgqFqymCQ+hStuM0kUgWmmjWQ+I3I7RGz0WW1Njcp
NernyrI4A+DFVp7hSlzBdJcfDpNBIuoALAzISaah7uVFUrklZOmKkvtf5/LJA7Gh
V8+0UvVXosndERE0u66A4br8N9DwH5y8a3D8JeNsN7o4Okok0hV7g/Oy7v8fKguu
qOUFkD0EfiEqOBUtlnuLVBCcNMX53bCgl4G9oHWLNmRGw4bQX7SNG5WchgXeXpty
xzyL0gTUwraUoG4sg0iUzF7KWCTZ/kNtNJlt9x9pWYEkWXNhENScWAXJlfT8dYoV
0B0eV+LS3kmAAlALdicsizsLWe+KXwSrpLhI7kA8dA7T64nLzu7VGjD7jeXOogoj
bybVE5B4wHJ9k6Tg9qC5BbQ4GYgLh7iYwpggJVz1uX0QZrk/g5b7wnQGR6PprYVR
pJ8kQd2Fmdj/NWIqRmcQf8U1Q9NKYBTJSMRtaUuy26Q/RWiKsifgki+WmV+SxEN5
bQPyTxyXh0nAAIOYMNZgIsZsYdCKiTHvgYDNSBL85RzeltARou9wQvHL/yNSEjGQ
+a5iu9vXZu3oNQVVvD6F8kThdgEL7tuDhYdsR8gbiXVI+gK8ey3XS/h6otfyHHhb
jcgURXvconZt5Je8aLVL7pbKn0pZHPi5fCKsCMbBmS0zryHNWvO3wB24gpO3JZnz
xPfGEr7pig0pLtKlepsG4O2TX7HSNc84tR5PACHn4tYmG5lnhLYZfPtVyv56JpSw
Yw3R3XOPt0qFvcIrHkG9z1Jio+J8rIydQfYqUH4Q6CXVq7WfK3mTb/W85X0r/iw7
b4nlyirDYG7vNTgXDXgChQFlNEfYQIziTx/Yme2lmL5I+kWpr8aOxLm46vtIyBwe
GWEt0e21E9UN/2suSDUXnpMTbwi6mcZVwUM7TQ1k4cMxJUUyerg3DkLwLBxwNV9S
B9/9m/v3yOGpX8GycuRi6CHM7l5tMbTyQSZKsN/FwGWuE3WmqysLmNYvVnUHZa8l
FbihLlCECUfAggs52W4ZlnWZNhEubhiDViLY2DosEJSoZJCTeUA1mVxZlyv7wq/z
Dzj7kdv5xP/eegjNEHFa1KoZcXCUGc6Cu5CrKE/1JRyqUxnNqcbJuQ9GyU/npcW3
yheZrrRqSWlcb+glxSslBNs0eQ5iBQkIfZaz+RSUxM2FORzxuOZV7dXKOuU+QPcO
W/8Sh1dUGzo4Pbmvcx4zeTSK80Boocu77xn9JvPg81/AkR6WSvriXWBlA17ZePb0
XBl3s2lMDVQc98N+YNC3h5FojYHBfq8TKGoxYo8nHd81wtrE7hyJQeIEEsPwVNa5
ek5n9waN3b7yoMWYcRo+RGqtBdjsAylGuRb68iLdNf8842pqkOuURq0GMdLW7dbd
+c/VeSk9OmNQmqPxY0wav7kBaMMqNjhLibbYOrhPCFz61uMdv7Qp8b2KNukmxKkW
w2Bk4wpQDxg+k7xyNxQVq65YIFO7blQg8lno4nc4Y8AMLMNobXABJvCsnczJKQuQ
taWHx7DIuVuF8ExqCC9dn6ca930kBHBNPoggs2E6V8dVBgog5FiZrfjXRGxn/ioQ
Fq9SU/nx4DYGKlYkS3m708n76XJjYBiu5EefyYGOM6RBe6a8mEBsn5JkSMuS9GIE
20RgVZAzG0oar93sPskN7SNEyBVHoEFR31BZh9gFEl5P+XGvD+PxJX76t2CiyTD+
5Ff1WiQTmi1bEQlijOEi+HWvqcRZmLMUH5aY/Pxji+LftJ61tRW6o8VTdfavHxpn
85jgqywCoG3TujLhgbn0YmS6E8Gc5TPuKMC2DDEDLXZ+BfaZhOS43i7jD4PYGr7w
8x7fwNKgD12/ff8jcMIh/kALamMNxgQE7NMjpfG1hmV0vWRyTle2QTcQmMFJ7coT
f/RppNyld+T2Cj8BgICttcc4iyGDeNa+JxntS4U5SQqSW7LLDQzleopy4bi5SI8H
/VT03gWGnjKM9qZuSu66xqab6zUnmlTR0hg0aliv0+jviIoJZsF+6njPNnk/pBSq
GBmDNuX1VH22OULLV9Hsikj6qul6ro+NKFndNDNiAB6aBjYo5oxxZrkQz/5M0aJQ
pa0Ej85vZCzoELRdJ017aMZueNO8f50hAOx0ooKwZttASbmiCx5MvVd/jMmf5TyM
xoFZQ+FK2xTqkaAfPpBf5og6dW/2MV+bIBQxStAsec7A09G93Cu4HeNRQdQpMd4G
WJHhUtMjR7oMFIWJU6uPTpRNfK5+19RifYQAwvYm0c4Svh/s8tlHjFe1QgBbeSum
1XirwFOblFAw9OudT0P7yfWAowZSRA/BMLc4cZTsUIGGRDizUxwKCnsEqIdowBPY
H+TuKRHUTni8/GWXXXJMojgWibFnI9k450JkQ6GwsUbeqM/TNk8RkBlvTNM07JgG
5me5P0DbpB3NNKFmG5aooHVkjopgVxArxGHw6t2zYa1fCa4XMhe6GOdTryvO0GV8
I9p6VU0xkdDLNdBJWO8GQy/alzVAqLyfADgzTs3JmuO+ZetIffjUmz/Uxr1P/mR8
oZ3Rjd9AINUpX+Lsx+TalDLNrAaC0foqXdgI0G3lyC4xlUlvouBOAvEt7h1SQLCD
oMpJURbXKqJIJz9hs2loLFQQZ9EnAsHSFP3ulpwB7neN+Md3roRiaExE9DJZ6ZDE
C6LC0KiEqJrm06P2TivNU+FUkxkvf2rewzCVL8bnYAN7brVqtTqmxYupkSF+FBx9
m58iZc2/d4jbhOeu6ecpk42LmbEOL+S9vR8/9SbF1RFpamAHCmxKmiKT5mBo/mKS
uBHepRew0s2jECc3vUnH4ETIWkInVlXqCprCMKwVazecvRV6WrEex1YabiwXgsiq
c+Mk44uRdMnSAuRhpkUX6GnCNMp61wA9dzNoaVNN3k+5+ZH0jwaiVWr0cwUO0Fkh
MtVq0cTSfQFBOQPIBqAg7NT5UTHDTl5ipAL0Gs0PMe6Mr78dpARCzvBXJ1CwX8o1
Lufc7Rsqd41H84wTUR7depbNVWuud2dz47aWVs4LSrAalgMa47bzYynTuqjadRUy
V/Zuu777GIC9LUfylNpeCUSMq+gFMWg3yuL7SvLAYn8qmoC77NqKNuB63A1TCcac
NERqj2pr38H8q6rA0v0WEAZB5IOKZTxTFd52/apf0FIH0Mi4ARtQLrVAgRPh33+V
pyuGvb8xMKCvSU3npT/8MQybDhpBjGr2UeaJD6Q33GVJx2fJyRw0JOfqByUU5jUQ
Ym/GNoRQc7Zzip+Ppb260FAKkrwBa4Jl3FvWJWRIozN+aJMPJhLEIFHe1AL4tE6O
l4b4OU0nyBMnjmbTEHeN10nQlHz8P6aNnaNigFWgDv9QHF+WvQj+I0nQHzEOBGhh
0PAPqkS8v5EVaVgcv2GS0Lsz84G+XpD5dWEHpKIDOoU1mMeSArEZGa984iDeDbHp
u+U1M1hWEdQUv/PL/oqdZFsxwitIaZZ5htP4zFqcgVrHSXVOrNE28+HMk1KFzR+S
+zQsyV5wTsqih1CPCE8B4H7C08+4cFCdb7O3Q9OohGXnvEOKI5zVGApEB1dNhed8
k+Ny+XywatTbA5Cr9F/bFTwat9Uyvmv8r1cFRNHf3mRyWM5rrp6zczS91KbG7Jex
dg/vmZFjOZiW1qkFyw5OlEkAE/PRsXj2FNQ2PRnU6Yd9vZTCHaTveJ2gOlozdVz8
5f/ivejHsYArCBJb54dHiLltivCdspcDrO2B15wZM50anG0agQ3VOdAI2HxQecrI
RP2HTX/2xozzHGgD2pmEJqZbA/D1AP/++9E1w0620U9RTFqFal9aDDe2TROoZoml
73wlQfG1PFPtTmEKUvrwDWQ7n+FIrBrHHT3piNOXaXHpo6ESrpj4M4ZEqaZ6TRfY
M8MmLzoYMz9eAwxX/Cm7WEts3BfJiWLtCFhkQ1GWqT+kBPGoexLizfkE3yeoHk/6
gPaLcPRaTKZ3gDPRc6g+FByjEP+jeSLotfvn41+DKGDKqXpUS6FYhr8S+lKlkBXI
NgXoIH2uivARcWKB6ivxdPa09WXpPJvaRKr91Cfc/Q96YJTchze8lplYLFbu9x8x
8krQpHDv6ogM4rIm+2pfp3qKulY6S4TTwoH605dCzA88dUKsvazjVIEiMIr+nlZa
Obc3Qf6IRGZOcCeYvpB3R1d57d2niDZTWvkuHZ026Imrh9qeHf9rjVXjk/1atvaR
xCO7mdJDAf8TOW/+CQjpWydlkgx9CFsPmHo/S2yX6gzRaW6orsaZfvMXKysYVp84
h4wmv+BCgqxF47tPCzBniZr9a42GQTwID54Udglt385Napbbe2u9vBIR63PdZ4lZ
NW/NfQK10n1rfnEjTGlFwTlHdBacV6/FW37IUtfl1Ndhi41Vh8XHL+giDrZ7W5Ny
vjk2TqjktHXAtolfbSU94sTWAEOSkIr/Fe6AagfbMx8axEltfZg8dzD7XlsAkpT9
KdRC8e12Qm4ej0Ab/33YtRaKk5bRnR5IMVS0Fjipp3ppAdsiQJvyv8kU6V13Ehij
GMGJeKGKzE2y+teJwQR9VqRoaDGLrYC6l9i3I2vIumPqANwF8xv6K3d2hbk8Qb1g
OrTnmKRAEWe/g5a/8B6zvywtgkDX3ZeiGsWUUBLS+0P56u2eEzxaS+AI9SUhsGds
kbGbSacrOp5XX/cmnxWop/mP8rCmYckIPTKvRAmfydPnRwNNcQaepS0dUQp0JlbE
S6altf0fHQRY3kTpadixOshLnC2zGNW+y9s5/Zb/4xwjd0imHaBKpAV2awrlE+6x
Cv9xDNr9DlINfABe/zdq/kGiokPDz4+DQ0lrhurX5AY9tW3SAT2zDCk+e9+XHKkS
u7QTa4h+/ijzwHAP0XuUIAzgnIOXlm9qBj2e7yAvJVT4F1sGvIZLwnFR3tVSKBDB
xSHkFZkP246J9zo3NMhCzphtdZoFaKeoDq15tHf2Yp0qpomJ0TliMdUpg9q+1zC+
ruBse9WKM0Bqeyyzx+aY9wrVZiTU5QJNGGeASxz9fwgX2nMHbA8jyYiEGQOXc3/k
VO24WsA/G1Raz3U1+1vUCi1d9qSdi3AIepAFlDhr9tnEngy9bH26tzrv7fBW4QFL
zeU7/evbwfXLYbhTuJVKxaIADpThF5V/Vy4es7ki1mpmG8eWVFLxQrs10EnZHE3w
9WB8lIpDfg1sF+Eh0ZFtMAHaUVe36a1lYB8/wk2MLKtNoq8QwSrvgfzulmJWx830
+VzRPKX+14p3jlqb1sF0VXvE03ghQb1tnrqKNdRP1Sk6v1e9D30827fcO7pF3GCV
3kce32F8tcJg8J3AMf8A7ienZHhIn93iMHq9xPgQ/AvwrHXyMXTGZLrXQoXIAUok
8J1h0glqplCBUxBhxG8EkmB+Sl37/1PIxiHFTjIXWSbTngUGSY0nRU5XcuHqg6Yt
tHdSvs6G3AQnc2RM7JHNYzdtbRKCvHfG8oJl2/TyUHTqUjXXwxomsNbNb+Mocp7N
5i3RXGPbLj+r32pnd7C9tY2h1OPQ0vLSGhHYNJBiYogFxRuVMlcEGySdNJjcx4FF
xp7QeX6zg4ZkNYnuN2Ll2ozxNLbp8UkyY34Na1nt7KDMmyZnRlgUEqhpaPQGtrHy
beP8VCy7GSXJnEGL6Q94dvcbhY2Jjrz+ihQC3LskBoquKbWZF+8z8k9OPjyVHpsZ
hYfWAlQfVACED9EmxH3cuL2CqibsGaz5C6cp9NQ2mWCcEzNM4pW4Yu70cacBung5
qbl+E+tz3qe9aRxIWEXVsAivuFmLGeNVysuRo/RUKfBV9EP3eonEtoyoXbXjS2X8
O8i6ZB6oqH6pKQYwYdPIhjOmL5lEk3TSJSXwqVZvlwQWGxbn6w0mp1llOTa8kr+k
wgURJAExuOUf4LXoeMWAyqgh6c5vyeUKBbGDQg44AU1Y+TUUqn4PJz2x6X114ASQ
hOCtVs9JWL/kYiKDTnE3PjPtmqhfBIP3s1lOI9v653flIb4d3DnIFm7Jo/KrQ0Mj
1s+ppR495hTlUNYnVPCw//wYrWXJTjxFusuw+BQf77kZKdcRZn6o0QOf6KU332n8
P9JlEsC7w7qaWWNV35WKXaGQ2aOyaG24V3pxigtqkaDqXYzCnp4eLCgyQuW9ymmV
KqkKjyGS6pyZD3MqVVjmkk51lH4z4Eqrs2VlviAQ5zqXn+S4v2GweK3VbGNfz3k1
786r6C6/kVRx/LCLOdLmnjenNzoaJXO2kLTvyPGF39QxysbUFkbB3MAed0SD7ZqC
Giypx1ju5YzQoNVkxE5PZHoUkiK+YfdYGae/gd4gshorU6w9ut3DCTSCcNExAnMe
2vy3j7BJrAdVvZo48BJskalsi+5wF2Ss0b7AZEOB8RxsPcUeLpBCjntfDrX7xRfr
bg3xpM1jsDVCYN0AY0EDlHtQYo/ogF4MfL69VtrBiWt3lyo9k+jhXQOlPiJmNiIS
uMAvW44y+0/txBLiXR1iDCmcqF749fF4Hl6zkyd7qnn0BInj9GlCy6MXZEXmv8I/
MznDxp4jvtiqvwHNcS0xU/jAao9cYTCr3NMeW7csXEbZSYiTw/OrI0EBkHV7O7/3
A7BDlDTe1KKJNtGL2aoWP3BpCiaK4yGne1Qem9BbXojxyMRxURnSSzp172UHivzm
7m8R6LMGDxKt9efcWTP+zqk5tbtcZBe0EnSyEOPzNpDDN1atP5BoAB+jQ9PBf2Ta
ihjaD8W277Trq+dA9xOfCBoFHD88D0kWnfUr58aGabACExQ5/oTscyLctnO4Xi6H
eR5PPW83ehD4dOuZ6YXOTZsx2sr/JiCecJBE083wrLBB1Am3pobpbqPIOKqOZKZO
biExLie7GkR2/L/CRI88+bUXWEm66osi06z5+yoMwbTO9+BYijn5jRF3CEiCGfw0
29hedY476XicfidzRFg0836wOq11T/9K5KRbuAV7umxhVNWZRGxW2sgRPVlYehHJ
Dq9rOri3XNcwDXiRoZRs9L8dVZ0QObVYpCl5PiGaYFVtEi0GOeElARWYmvQ2dXGZ
AmJQEXaJMkQoTVAqPKUdVvdkDlfUD154EkLBkYdBd6kUrUHsyEwUJRVQKJr4R5t4
etWWSGtWFP/pskAO0fAk+0kMmoj0Y5q0NR9IUvQeVtrb7VykVAdggZ0LE7o9fv73
jh+GwFX5oFvNSLxyjBQwEvYn1ATINJ+c/cNbQOeGeGeNY2NJtWSvBkKLxHjrJUC/
B2KiGj0iRtkUOYu8wIKFUK9Zfa14a5vfs+S9utpTqMTxVrq9NE/fVz7rAjvpWtiC
/XZV/LZSVNXhkkqcUe7TK2efNtS1IV+OcvHEoD7w4eDMm9zivBe+rHW654LAhUP6
zhcF4YXX2Y9Nx6cTDpAzNkKcoNyp6QzRx6NqEkR17FmRwLy7p+rcJUinRLKDhatZ
r39rwpocfADqHTXY6qZsAFpUkaYQlpGAk6pMILluS2kY9gk+WPrTWEYQZsWZZHu7
opX5NVL9FBIYrlMFUoIi4Vt37Y2ICwVGnt1NvrdN0h2xf0BOXkMWI0N/JRISAWl6
BI4l8qs6YaFdeq+rF0EA38CElxn6JdZ9wnDlokthoL6hUYknMCWI7cA8Z9drDNWY
ZcwxezbFsbn0vKVYehQBEGasYHkqjxxkOZDLNpIlxUS9BmbTerVn/jGqEH29ppYL
jyIwXDK7L2FgV+Q3kWjdfF/kt8jIb8V5WptRQfWVZpVsvpn6ymYzmrHI58KO5uNh
iHaVtk1BrkYE5rydvSyhjbK3jwDTN13cP+Ak8lnEsQExjTrGU7O6q8kgmWIZhiXx
sKZlKbrxuXDTg5akNxmSrAov+HMgA8U4qvBjKq7MDi0s6iyI6tQ3Deg3Abm8FLxU
8wxCGU7NJ/BXtWv/hc00ZawWskjURtXe3EYYjUh00EQoZCm35waCfl03QPi9XSD+
Gp64LbYCUFub0YDIB7oH2nlPGAoU0v5uumXH3WP1/SFSTIgohsjoAOjCArLd9pjT
MeTAC5COdOYv9bV8YgWI1JlpHfq2ls3hCY408K3cnSp8d8RFmN5u5Z7otyX2pM6Q
oyS78H+FFesmVsr9WPikA2f8jK+adYbHEgzJadte4nQhSLVUSDk+HQtUQzRGI+sA
qmob6Vdsh0Y1nuuGpoAi+ZQDb/P3BS/cs26/kUq3PMNLo2xmAu9Z1nD/sbnRj6oN
4jUELTrhcB/kAU5ZnxDb7KrMvb2TgHjxGSmPuluI8kqir84Ko+5vMKsKxeTpTp7L
x1yGNeddljyyK3LzVjFWqbfLC/2ZRRRxsQT0p8xHdQIMNbxQAkPcNqsKenev7HqI
esPZtfZI5SKwGmIf9boeDN6dLYgGeggYnRrg+WVi4BESw0OiVj26hEn35a6ojeGY
komG7uWYFOirjXXwI3IJlxop7w7hsTK/wi494OOJjzWaenRRxoPvJ4tIUDIv7b+P
32H+y/gfp7FfkjwUsEgyvMikBvqxfmFFbOSEn+s0joa6uYbPF57APVXY8/rAfo6t
0zU75+HSwwCxS4EA+v/A8LHumrD8IX9Su/UeMk4kmdJcuEIXzHyov8g8HsyK69tg
TVb7hJiPz8JQEQa41WbAVH2dtDAjegpFvtOPgLBt3rSRiQ20bPOZfL3HxaQccw9X
xvUs5njYr5vVyqdiEHO1GN9k1SlYrxh+1S9PKR1Do4CWPKep2GLdqx5EEtftmfmY
kbsqzWLGtTbzgmL8pO5MtQRMAxRQuXxHF5r/ueU4fsZQNh0sK43rCJzYJG0K1QXC
auiEYzJI3At70aSgAZ/opb2aVhtPU2gZaarMgxpG+iq2TxoAv96V44gf+YwQDIyW
V6rGKom2WUZDl0YjDBDlcGY8cbSHVPUMgAgZo7OTvdfmvmrVs3dMm2Q2xbM9PTNZ
WghPQQ5otKJQLs98NhruSxEmMPIuJG1m7RCpvWPswRsjpDqa75e/vd8pPbkJt9QZ
6RQBgOLf8hvYp5s964VRCTKtby2fDP2KQfBnCpevqPAhmbj0/I2jD9Re4WddHEU3
uCzqLB3Q6L6Da1oAOCb7bkWux5MZuPr1WKCaWLLta42qMQLkXNQzNtqNjf+nnVm1
rJK5ZfBEFX5C2MGsOQswry7sl5kXfXb8aay8liWIxqc1Qaq4QM9iCvjwCOf9kunr
qTS3aB68V11/U4n4imr0iipYWh1l2c1x3mixaEQ1xn0PscnbNL/ulf7bgZjxe4Jr
qPvCmvX0xePUmUuCVmx4PqozWIzE9cEarBbnAa/qgGYon0RUN4gncrxhRa/t+kcA
n4d0YNLdtyUiQfqbG4rT+zI1phwuLKlwld3LqTPhxNNTB3nck7FBiuvMgDFxVRgR
mSHLlZgHeylWmAahP9JySr56BDJFldDhpS5BhsUhYEjkGILH5rR++L8CNYN4k3Br
7aCOjkjyXUyOkX1itFZJhaDIke/hQ+bOTDZDACRAzH6e7bUe5AmQFetT3fDinx3Y
OY5RQjWmg6GVnHdYXQXq4EOOBOqy3Ja88X+cn8Coz1ixwYklBzo2ASfRpCORo4sY
JPFou60x1PajbF28ptkZcwfFHneG2ZTWNcIS0OhOv2T6Fe35IwUrRqpUai/M/19v
OFSBYWa+rKyKApdm/gA21pANrmPtTrey78fKWqba5/qFkueJnXpBGwRKqDyD1Hxn
5j1wKqtDBCmRfTx5/lKo3Ck9hQKyD2IlLAbnEzNeeswKezSkZ1t3W99WVgiJBQM0
53rHJHOlq5n0pxKcecZw7w8BNZIIUXUL/axlswYMdeeGm+BXC/4qJX7Wt1IQF8Uh
3pz12NidSNeydMj4n7bDxv40KbafMxsdrzU/r+G7k+stla2UTpYDlRw+vgfQkjg0
7CJemXuXNT079mRVove7QXqu0u0+cIIdZ8roLVTOMtzco4yWNiFnGhDV7S9BgO5Q
yAQ43WOVY2KCrQ3MHZ4d/v33Wx0iRyMEfnHMByhfNQ36dZqmYeJLzaWS6IGtR9aG
xRcBCGa8rTg6JQ1fFKeK/N3iV/BtJETUiSOa736g5ieQzvRSlqRUv5XUdBOTt6Sj
JR8Cr7fEXG0V4Yyr8YrjIcy63q13pCljeYYDhqluJ283srwdQL8vJ8Lg0JjrWyqs
+JfIFYsUZNOEcamHJH5VnPmcgpvDvuQe1jQZJorLXmhGjpQEBEf1atlf6Q8kwh29
qRTjKE7a9GG5cTrwglTMBcTP3Bs+m9reQ3fScJJbsv6CF22eY7Tzvq/i5u8ho3vt
CJ4OceA0fPWHYyT+RCMQHoC+6TszGit+uw43GtLTxbyLvfI6li0U+3lIyR2zDD2T
B4afVSkSpKyr9JJbw4jZRQl+h/aVDEOGKIye8ikd8znL1UdRnB/RosUFtPLHWwZ6
9hFwShHTjibRAP7jqa2TwqlSPjxvFybrFQ8ZJJaGcQKTm6TR5yFOqs1K26sWS0fJ
2f0ymRudXNhomXNOpcGqJ7rQC0QsO6EgpPKSvY17SQCaX+/8+U36mGm7GlkE+AOg
OWrYDGj43otBeX2sirgDyFY1nYCBQjdPB5enOp18KgiV6TIezBuHa62Ka5JPmvPy
kkZSRDyaUog0/Q8OZf43zBff/HSTi91oZFSKiRZOwYJGxO/LBkkjmAcrWrpK7z5H
EX1OndbKdlvMxQt9PUeAWeFiBEmANhmqeD321mueevkfuwz8nu0ZSlqarwCIlP9M
z0Pk2XKqXVP5ott8TZgyNn4vgXTjZ6ctDMUDpqKhDsxUeVwj6dB/8ztAP9FXTBek
UbptagZ50E3v7a2yFijNp1rRV8GN1c0l64Ae0oj5q1a6cgp7Qi0VUxEYsFrA0Nlo
Qs5/N/obi/VBFTI/cGERH6AfENd3R2Zp+53cbkiE969hUotDtI3VjtlwJPEgQn0S
DrgH1oT8dxVzSrSkIB+O8kL+0PgApg6l+fzJbMtSnjuubX3z7Xx5IrSTLiS+udPh
cr7NGmYHLO9L8pRiHgjiF5FaEva63l3MoPow0TP9pyOapnIa33omWR/S1ecQqdEu
rA9ItsGF7zEzlHvw54N+mO9oHGs+46+hPeGYllvlgJHHlCLhhN8hfUWHtTcaDODM
w9TRVx8iIW1kmCq/EaJXl9dKkfY2ahVSNtEbyYEI9oP7GANKK/CxmajE9k04U0uI
gO4W2sT1IuqOI2k3IHLQknzFKq2aSJZ3/gaJbIZ0PUCSbPby1kY4EdItP6SG8eID
n7GzqVIZ4l5enHyXQOx0SXQTsl3VavE+SHz756AFRPFSraWK021VPJndcmb2E+XZ
YwLXktVmMWPccD2oHUJ2xFfSQvnEnqjZ3hlGRstW0FenVHUzRLFBxwQ7KZ6j60Bj
KvWx8MXhMv7GhPWkiZ5QrImyTMN5FWj6IXG8x04rxKQNNpo7Jf8CUqq2YM8gGNFf
fo7snX5Wn4kVZPk+hhR26pj0FGoJFPOlF7qZ/y0AGcU3aBvyv3+rME3SQ7LU+9qn
a2LWq+bhYtFKSJYy+r17jsxr4JQUCs59qRQC9ks8AnuY1gMYS/tdLtHB43vgAHf0
qst+pVQC2LgwMpx+xzVmS65R8oT0vBJ6Rqm22a/3sPt5Nm6gixlkK1jNBBxGKbKl
jPXQkVY0ZZu3B+9QXRxvIfikimi49kK+jBrnNGhsOcmbaze1TgUzgwXLphOUnb+J
25LMgYv78Rvy96Dw8QmqsFhQyLJmU4HmZnquBUxUblxMrm5tR3zSCvUSr69YmgNC
l1avOTVtXyDLLn+aeaSzZC269tkXvg3jNyAc4dL4syqg/BP4PpjXJLfBSVSChK1h
W0CHcbumqKKv2Duute1LenHQUPdQsm40qyv3SFZB99RMllote/qEekwaKmNKO9ZB
6CMSxd0IrJ7yaH2OG3TupKTfF+w4ss0lIyYAlRjU0bPrNNQ38LSIkm/WHQx8uty9
xK3q29HZWrqQMfRXQ5DmlO/krOOMeN4RXmuYQlN0LA0SxV4WKJf/Itgai1D+kVqt
EcPeu7gltZ5Xm68gyhfpSnxCCHv4WdqN9/amjdGQt0EUNrD1LpzjXlBa0JHhi4ge
DNFbZTdebqE7YyXeO5sRWPInEO8mtZtLIZep4rdDusjmAwVo+xqpOnw3A0DsKi47
EAP35JvtWpcKtyLKLtQzIqBSgy48vPaqPRXAhr06q/zeM25gZ+iTZ9KloIDjD2RI
YzavAX9MZ9zrrahKdNP8hr9jj3FgiQPq3YqgkNNKxxzFerycUSFtVy4BSXhl5Ci+
rQptaSSoh7L1to+K/odcuCQ3NvGrMTwknZfa3tnGDotbudxApqr0OBdzlb0Qj83O
WTAplMpq9R6lGHoMencKCMlhGz/GkBNIZB5vzfDA8+r8gPXC+aU0PtIDCobwEKsh
FA++lOpatCEUBqEE1ZF8imdyNrBjwLQ9d7Kl/Nfj6MVBS2VEOwRCJ7z6ZqMEhSgp
LKPqhGuYbRooACAtC4j50978HXGrz6pSOdZTJd4zc/5/vIEeoltqLUm6NrIjNGbb
Ezsr1LjOjBakhKTDMFCns+8bFngZeSwn5q9bFnjPr1CBMPNuOoRy5JfL2V6qDzPi
CJ2yoE82TrcVYovKlyBeKo2XK8BWn6Mp4ShiWRBfHcocJD0ImDrh0yYqfTEse82i
pqKwxsKivG8F57/72SSgH7P7NW8yt22DRtOGiGvXhjostGVw5Q6sioPpVveYQm3I
5lOG/J5peoj0mAwTIpRmwyXdySFIACPnx7nFxSRxxPKs4pNsHBXux7kCV7jErmiq
UTGr/+v0/NGldzQUUL+WSYQTDYns/5YBdx3+UwFClE4bOAX1LfQIUudB/jfmdCrl
LvCyx+t1VTDCfB3ibn/DivAGKLJ7GVd6qINI/QNPDh9kfgYmoGaCWzgjY1PXAeXn
ksSPIf24y/pYDCdfhRCGuucyoxnbFoq8sjYSBPAYWyJnQxlsSQIm6NqtOBjRV2tf
kkYx4l5/YRT505ype6b4F7XHH3AbkNqVa4h6PjzhuSSlQVmcMKBJcVJA2fA9PH+m
2VFvrht+05s6wJlb0cD2v/q1+UGXIe6m/jcXxJMJ06pldvfMdKVtTHlHNSaG0niJ
PnK4JaFIirvVnqT/qejDVH2PC+k5MM60fTBAdGNXXWi70ndsN9QGG8IASNaQET+6
FucCUCuJ19/+icqsfsgvj/rCSlhFMJNAjthGP8/YLggxu5GBABjoK/tXlFUw/MP5
2w+aG0JeRiqLtt6UQevJkR/y3Qy044hQTS+gi0dOta8ShbHJhsocQT57NFJ2ljgX
XDDEHE0L2tYu450VKE02PT90dYIh4ZKu6RsrBm0Q2Va2HVVLXh1rJUWNVtLja5K7
T7eu30Odj2LRYEG+011gjuix2k3LcvhBV6HPS8q44WK/kS/jHsD0TKEKAH+MHIdJ
ZC28438k1EwJsDWY4/WWnf3i4QeKVzd8T3K7IjlUssZH26iyrZU6Ncd7jnOmv99T
slbDIsJzxRl4qbfG1fHiMb6Xra+y4uEXj21dMTjfqq/5RtXGaACTZIh1etdJJMrg
WWgIpS94eC438UxB36KPci6Vb7K4tEt7EXX0lOOsranpiXdHETzF+vgdTeW7txCt
iOjiSqnwYtIkCAdr/MQS1ewcHuGg5XVtcr3xzCH3zM69EF9OuzGdLxYP1dlriBX4
hn7aTxQuCIwzS76mvTq212fev/S2QX/Sw83hc+0BY3MJk6TbktWwT/rbgWIkEG3c
hPU8IphoGOk0ew164T7MfIUdNibCb/ifyc+GOcoFrhX28p2//HJhMY12mL2UItJ6
JgxQet4qWprK+3cByJNj3IQ6m0eQMs1zAkckVdaeWh9qaD8EV6KX2Qgpwwqf5XTC
NWZUk5l26Xntx3PXqPvLhENtayfL0nZ3w1izFi1YfyEBA0ZzNPgWhxQ51LfqTUZZ
KYLPBS2LE3qAFmq25OBlXqNfs9sZJGqILdx3U9bAS/COQU0AJVPvAQFsDXYXdrT7
zqrMNxyWhtJYwfBKovAjeMWIM4c9GPzmPNDBxSNQHECcKC5m0X2MkFf3qpC+JhXf
cge3zFbdmKJ+U8PZYReBPVS1gkw/hCzxCSnn4w/4GMFQ3dmYUBxR8fU/MXXV0Bcb
NQAeIrzgQY+cGAp8/cDrOClFBgl3A8e/1AROp139J8EJzCJURLKh4f42lUeOnUWL
w1drsH3QYR7BGIbCsilF+b/TIQiweO92raYqefwVbkRtpjw7IIx1JeO/PuwRSyQ5
aJ9ySEOTRMxLisY7cHhKHDCW4MDVMmUtDHkF84/iCwL0xgyfMXGa5XVZ0pqqcibm
ZqL4tadCPvwyC48kEs2FLXZS+BNOifHhsCkHxgRwz3z5/JiumAa/N8L4Yo8/FPBw
2Cv0qpulwQ9FYE9j/wxG3HlkknQf4pRW8cErgH58FgEOsPUhchBW+1U6FSpvuJ/Q
3RBDydy/CRlH6A75tve2qB1ijYjsVMUQpM6OGHj+KALWAmO2ajL6fvzHMqqFKJtK
ltXQLLFd6KPYWXdQRoTNl0SX8ukqt7vmZP0lBU/xbqoKtlxw8J3GMqtjDRtmtC0w
xyHuLOiHgcGevgsq/zAIaPL3KQfjZaBoE09KjvvZpKCgueGnw2gIym5fve7UFJx8
04UtA7qroyxzZeEt0/qqY8G92xUcqawdGDUNT52FH3IyQej0uKcxpC/yT3IR3TQQ
3St8Khyz0dWexVDivFg8DYWTgxjtaY7uaqYotp7zU/0cqi5S/Pwb1haUxYMzGF2w
if/dyYT/K6TqEE1dpLOopAtfRyuw9QWRqKC47xFkWmGZra0zga+P5bplnWwLCgbi
b6vHneRDxBHcJLc48ZzYxa1axO4G72SaOwMno9nL7QOasdMP+Qo7YZLr7LSaRbxx
t2rROrd+ysh8ZGrX/8zOHTaBwk6l1x+cMYFX5VWihYw2Gze5vV7Heswd+wzCb7Gu
ootpZd7PHsMngwM2AnKBHDAA0QVQoFM1n66HXB48XtCS4btUyXEj7w4Rc2ksqWKV
6QDY+bavrTyy890j8MO6/zTLjHUkVU/4t1l84+sJzGObYOBu+wpOsGwZzmp0A76k
vW1ZSzgzzWoFBJh+v6g5EnymspZGB3fg05BlRwlqkeICLmommns1z2oy73hy6l9Q
Cx8HeA87yRaXUAhvq0OCUnckbi1GH8T8OmaJd1nIuS8FGEfhBObkk1hZ0i37ZExN
QHkaDUx8MvuysSTAxGHDzlwaNIns9Ev6ytu2y2BpTJocUEiUyn+eaWrwxjS8l4H5
RqPfonUkBDelh/2GRR7AGF5IK4r66RXYFvxQCxOEbY8Hd4X5mzc9g0v3lLicZVN+
lXZ8RxoPz2h60iF6QavvjJMgE1VFaI/s7L26sKwVtit+ZSbxDcOD0NB3cfNoJWq/
RgprFpDS3AZlebmXU3iZsoKx5vcxy22g53zfSDspQEvYLzIzvTLO4aUyxUwdYglj
zeTc8opdQlMCMKPtSe6mGZO9GsxhTrSFO7HOx+qmn7Z3CTkUfUgubp+2jhZK3aPA
hB3xwEp7bda+u9E848fFtoch94fYI52ax9dDjCIUmfBC4fyDiCDo5AuBAgeiNt/b
d5S35qRLe7tfN6fQ8B7kQOq2ai7fOnPzXHmKXyQsg0jFc4fkow6/NfyLHOuL6v2i
IKW/yy5Ruqij6lzXUCXhHqUPef6x9yY8FluJ1SZmr+wVY2PiQ+e+QgTNN7ixlPUK
RaLTrdFyhHRhWkWdJ9LKRdyG4nxUz6QIaoNp+tMo/X5tmBOwbK8ckUaEVGrYGKCm
VPaxN9t0EdWiTZ6+EsLZpI6g5C47DV+gi6aSQefuXB16BYLilQwpTDBB5ONtMfpC
CmXRoRy8HsGGydQtUuiGy+EKfTCCnj56E1DkmN4N2hMSeuKz+IwyrJoJxCviMQ7a
8iTvV34DC2/I2s+nPPCnRW3G8nuC+mO+zVnBrfO7t+n23mZ69WVGCkhyW4pGt5tD
3Wp3WkHBJT5GppOQ7R7kz1J5iJbCIQ6xDzyEOmGWh04arB0iRB1MStX763xWIAte
j6WSoUAdVXkeyuENsAB6USYXb9pMjHfVDwCvaZf0lD46JZIvV/aipW0tgJwxVk0v
+oFpWQRsxW1BGfGCXX7oskBpZnB4LIHecypS6QWMijBdTI2ZlqjO0mG64aGYZRSF
7ZUwzug9nDw9V2FkBjyNmDUkqfS6uOU9cvxliM4CaxFesKVnAmowUi7drkmuQGew
TL8evM6WUKSWDPVvmHmcG3SJZWWDrN2hsQlCnlucx4wZsqh1eIPTov8S4gl8LnxQ
4T9QPZiQnSMgOE/49DtGnn7KPjqqs+7Mb0qpfpQKjQ7pqXxs7F9es1+cwBPOTRQH
UVk5o0hlyQOWOPh0qbAwhsrCclFQxKghq6B+lHM4h11OfDlyTzQBjdDgGcXZEC7q
8JeHfUZlM+OIzGECU7AdkwngLdS9BeR5Wemuo4XkdQzYN7mbScgB65ZJX+zbNwDq
l4Kz2tPRkzPLrE1Sk9KGQNsF6fb7/voEuHAdjRfEdk2VCYplYcEbRGmHh1ypvp3T
k/9f2oyooZotcsVE4VkHIqMkcWVZThGYckSzWQgaXK17kkQUjnO5CSo6HzZkTpun
rklqFQwx9AYF2xIP2xbi69qMLrckSxgHBuauTKyT8ESW4naTpPzzaL3oL5kSX5yp
5Uf+DEYO2c8ucoMQNM5/vDdW0W50isbztbaTWh5dcrE/xVC8+4d8E1cAnEl1x3u7
L0HEbzcZbvcCqZs55THlP+waWLWNOr+5dGknoQ4fT1xoIs6qajxmotAjWXwwMgT7
updFqCleqbskXuQ0HQ8E0RSdxUaWAC/13n7GNOIbjkypbQsjBeMVbhqFG7ufDdPh
yd+YP+HbBeC3CRgFyHpvu9IOvO7/AgRNgaU/hfeGWqNFv+sxBfZwfBfyd0cYjDs4
FAYasnVnzGBjAd9SN5MbSeDKD15en22Q/EKwOmBdfR2STwQ8aavySm4R40Fu6kES
WrdwMXs+0JbQkbUzxpKgONU9A2V76raVgPhrVwN+uOm4ywdCho+pkjUZNbi8ciul
0AgEcPbnAlDpi5LKm8MHgULtRHCRl9VFpk6+cfGnHXI4PfHwOGdxarFOjMF98E0V
5OG4atYLsI++il4NECzMfIXJcWHUWZnCCxYMrtGRgHDWKMOesy1o4AbmMNnDRhKR
CfjzeU7pqfW3laZ2G2KjL6jvfjAQVc/k3LrV5Bve5kd9pv3NK/ZwyLXziapo8FAm
A+YW+D6aF5oTTH/2Yk4Vzv5uCICvGnWyxrgry/TM+cQqo4GxgyB608AxRBLkxK0w
yYTUn4TxhXxkM6eQkir9Y8NMwo6HZ+jLSmzyQ/8k+d5PyBTwY9Ug8GYWldNkwVxh
JQYlnwkq1buhNy+pjemlKZCogX/Ni7PR4uI8E0EanL5BmqPDoGW47KwFStg4DbBp
+l5g4j+UP14OFpYdO8iZnPvzC7UkJ2Oi3tpiARjrFp5EkNHIpXCzLnDLA+igqTAn
/pkyJxEt6XZm6cMpTXgqSXbma6DHvebhOr4viDPXNcdO/6l7DcbKJnjllTzVccji
2qi9htd0pXfufg9UEVB3vps9BpLwo3zoFuPlYCFPTIa+1sp6hLLnuJJq0yD0oc/U
FpCRJKWPoP/uWRHXYOiUIN1W2d5S+5E2A8QnMEVEPzLerN9QPAJi2D2zQqPxrcZR
PIbBBN+Dnm5tCLy1c4xio/H9McTFSlrin4Uc8CxIFgEA2P1sB5WBf1H+O3dfjoW7
jGBbxv3TykllY7GNUVL5MYtCTvbKnT1Jo8BlB8clsdJINP9ekoGYvF/WjWFkv6Tc
lWoCq1jLZNin1eMbqPTNAILauW4zho717U9ftANGOpLNMjI4RwPCEUZ7mrG4wIY8
nufG8wAVBsTh7ZAwZcdeIu8v66SdsyJc8vcM4jKJBxDFX2iDvYrHN1rdXn5rnWVb
/cWPdPsfnzsPHu69RfeCRVNzWa6b44EU8YR7ks0HnSkRW7Jkcysncm8WGwNYmh4L
MVqpYs3wp8WCtAncz0t4H7Lz36Q5YwTndYtRkeBUfF/Pj8SJVD6sBXtnG2LVzD0+
MdH3fQpsYKw9TmXPNt7KRldzEWGKZ85ZXodIgIjoJjdU4NSHOhvR2MXvi1pozcnc
FUwYGKc8rcrh3BLury2Mpk5GFCPCg4I4OEd6SQM6ar3uW+WXxvx/oNJCCNneje1C
o+1QJSXqhU6fu6dGM6OlXYvWXcTj2yDa/KiiqDvTIZm0BVUYxo+bNBuD0FwUEM6s
OFAOxWFr9FG5LQBU2KPdesUxWq969pUI6CwbhfDSLktdz4w8ceXRBTt6XT2Co/TI
y8TIraxbvyMnu1XYTVTOkSkUdlzLDy6RMK0sgYBSbIbYes747i0SDOvKDN8c9Q0q
TwEc5OEm/IWBufIKkGLy33VDO6rFrwzbuQtjdAaMSRDYadUkTnsMkeHKMpnE74eP
URyQMpMc9/y2KvovOC8WYYedSKmTQB/EzvPEAouX59ooR5pR5vrcyq5n7cMD5TF+
dEluMdZUyhby+k6KuVLd5lGIdWdN0I6KL/1JJS722kyGMhNJaslqruulQ5UtaXve
nNSmEvKFlU6yF8yvE4Aft4F29lla7uIu5tzlE//hDEL9wIPpoNs45CYLOtnhBU5c
gkFvNGTe9dHQym8v+o6Fkw5kxXwAtGxlbGRFTxo6Bk45D2EiVn6DNuV9y3jl4VHp
MCYuioU5WeiTQ3TF53PtKTNrdgv2k0xkM+DjZ2pRRaWd8qCiLysiCWDZEFRHmB72
OPTFzo2xqBTAJYGnb7Wx52zTJn6dM+Dr2QNlX6RJsl/WjyIUV+QgrLMl4YjTE1XJ
h8PKb1lLthtiZU79XnB21xAhIPLDvr0oVIRtiaJp0MekSMgWnXX8FwkfWcO7GE+6
Yo/e8b5/+6idMFPq5OmF7DRUnsiTCBUGbYgIQQ74BDcndYoBDSHQOoSz9KjSOoBC
pS4RoEBoUTnB/PJNzw69mKIYkbYeb/yIwwFGwGiqybF0KOUqDrIHbiQUikdVg0Ji
qAwBtRMxn/TwUJOGxOnuYEFDIeVXOpoZJepYbNJv92bxwwzCwjvsDJ3vaqvJ72l7
LE6y3h5k+W5YdnwtOJZMvVEyilOEohKp2ChxOkjirIA0zBmfHTCJfBmFEuR2B+Bl
z0zq9yQw4tukJcNbxhTgxlXEoDMNwAS4rGbIg2abZonjTulO29Di8L1pt9E1nO2i
HOUAd7MqcEz4YSU7hjA/OpalsAcFxW3g69QnBAgG172+zjf8ou80h8+PS4g8nobE
Joky9AThxzIqjw+ighjfFcfCnpCS++mpcvb+aYxPx9bR+kvNKCtOFIDXHeuiask6
DOZHzmElO54gjKl0D0GFpCN9C8jvAmmTwVSAAF+Ps6/WSsAr15rC1CmbPmC8fOWU
Rb6MOVlEZaMwOj4+mVrBIfZqwMaBN0HQw8ie/wuSgSUe7VG1b9wfFRdwiHBKIRRp
C/PRx5hsfCQZRsMeevBLJLmMMKKHA5mwWiBGlchYmfkHjsDqs9hNih4nrn3ac0Cc
Gb4gE8DlQgPs+UcQiLFux1MoB/Rg2DvkqHf42NVT9hZiVBznJiAjhhcT8UqSPJOz
I+W7rvkmEvQUArlK/WLrb9XAccj1uUTLtVGh0b6MQPYrfRQEoKLx9hDmtyPR/k+o
JunyqIPg3N6G7Mw7W67pcaobEPfEXCTzGqNfp6EnbXc9pkeQ5dQQ/BQCaA6P8N1N
660jFln/3btkCVc9fhaA3uCIo+yHaPPXvYHMw7wtC4g35L5UpXXTNPHKbhp68GyB
8dUVQqwpeh6VI0kjNldHCakt4JAf/aEWR2RljLF3PLObNKXSz5yg+QaLhFgTC5fT
0gWselzteweG+jjsJ2zMgAbv+4j6qXc3tY1pnmzKHjDEDrdkruHMfUxQoBgflss9
HkgSxEhRqyLXuu18cGlXaQTUJzIuklw2ZBfaCZN3wsc361NHi7mn3R1Tmp75f2R9
Gopgq/cy8llcWfVck72uh1DnBZQ9BU4aoGHpKZT/+txmNHZDdWDjMMRPyu5yExm0
ebuzRwxxx2cQeaoy6BALL5Nakkwj1orXQp9vL5ryB8ba58CCYJ8+T1bk1T5zsCrL
wKjABAWTFVQAyrvsEJ3WPZm4r1vp9FBe8w7wdpPa+XZ6dFv1cbhj4SOhsHXCBUkA
DR+J6pQNWEbleZbYm3dXi8s9Esb3As4oo51Io/EQTsvC8N6OpdmqR3xAVdDjS45z
oipuu/sy44NpRHDJmT/z9GetJ/5YSEA8pfXndPPVpQrifZEoid/2YUIeSOpaJOv9
1MtOay1rA0Pk44zzRQk7AXQQCJakCQHBuDkjgDG9Zrlw4GrdTZ1igKq3BHaj85RT
OQUfSMgfvWDHOndQ4jlUP46GPxtepcGqeYIO3FbTt2rRXKWfLvjyglMsuW+s7+cL
hF7SN9arnSVs7VgPq0RI/UyS+9s6IPMPWuK3sRCJHfQLQVX8QMpiBuEGSKwHCHhN
OiQXag39t7AVWe2fA3l6V7bOUJynccYJCvDNCZTOtnPCINQj1f3u2iL6qoDESSw3
gCw7FBys0idXBfPNiea4t07enHM+0Vvbd56HTbL5JflkSZf+YmumI+vcGucZltAU
u4UcmCi+bS3kjU6ocL52tYUNfO8HOicrVEwzWLZT31rEaWGc9rFIazxD9Zqc9zTn
fDdEtdjzfYkEJSIOh3nNMJedpnEhUS4+js76Qmb0Pko6DQVl9FlCzgaCtOHQO6c3
r03K4Ta/QSnEJGKB8QXz7RwoPSRKWPRkQZfDUySOA5iZWz1TzYJ1NnU5SpefmF/Q
PfYceqA2mvUsDzyijExmKVA8WuJNwlbAPhZ0rSYYx6teUpt3FKUOCoGizSJYfzmm
QnLaNDblKfGYFbfRNoxc2+JJ5K8HlJ3RS+s3UavcAwb6WU5oT6DQJoaOudGRWtTk
LR+Se2mtuUn3zTm36hvDjKAWfbeYOa3zxSSoefzkvTyYtbs0VXBa76kmkDHhQnHl
gxeK9zoongATZYWZx+kvuo3KCdfQDpLV9hRspeuLknB1f75/PE6ltjGH+chC5aUm
LOzi++FewgbJJmxbEGoNvTbD+veKB/h0MdONHOxh7PDt454CB9YyHFVTBVm651Gr
LSROcLKpZDtCvcPX8UfIZhSMaMWT+hkghLJGQOHEiCh8lxTJ+EJO8kkaZWXbRlgV
naBPRQYCBvE9fJaUe7lpewCbMMsFxj6VpvFoH3uZmcv1zzVhlBAMJL+EjbL9GtoD
LG/QBOnZLDeTYQhFVeEvekxsKdGB1potjmz9tUoSvQF2w7FxUvSGZGzzBi5LyTcG
LS0HDCE/BrteakvMmQm08uUNXIe/vs2rktZ5fbEwoyVPsE97WjZZ9pK6tZSDI9/i
+rmHNug1mzuZccccqFouJaDlLwvltBmxRQUPT+SzRDFJrW4sg0t/oGEuVDUVv+3r
HZ+GlN3AydKSiLyGhcT316tD0SQQ/9Bh4MC8aTnUm5e++7rww6K1/7IZTnWwvmbV
ZA80XxBM+ylC0Dqc4HBc0nt64tBuj38q7nbP6by5i3oqj3BgzfKKIgQdVd8FVCVg
9nynm74WKxbeXB7s8L8WmSyIhWg1FPDUwtvuqjKyF9Lj0vWoMVScsHn7CQXMKc/r
PMcwNPhTrFMdJVcCbbBB4iUbeqOUAWu+0bOoM49g4v6nSbBO0mYESewco1u1oT1Q
ObdRhZgZxB4lRULauWvHHIl7EhSpTJp3u0ALtwZLLQ4YIDFBAQWInR1R3ssusaZs
m3f4E6HIqIAsEY31s0CzXe3zJ4ostdpQtKQ11MmuC3txdUqhkb+yFDqPKOC8G5+N
qGvbghFVc7efySgetn+tboBmjTM9pyaXgsGhMshWyOKajpQDTGMRQmoKc9OWcfbq
7a6Et69SQFcOXpY0HlhdtnZ9C9XGbCDzKgGS3lRX0agUBc2REaFp3r2YrjOFJK2n
FC7XywQnwsW6q28Eadlcd+OzBwNC3rpkqRZsdbQ1F7htkcpWqE0BRtyHUIEcE7Ab
XvHBkWlTPy9irB6+Ru8GcQVaSGrFEnVa3U8RoOzr0fCeNrY2l0RSw3jo36ix9uR8
TI4JbHJ+spKS07d/4VJ0WTs0Kh5bl4r4CAmlsvD646b3VN/ISFe/EqpDsX3v2GF1
732mHM34hnychMJfNsBogEh3P0YBNMWKDdYP4JwgRfA+QDomTJdxPWoqGsMZNLUd
x+z8KCcUvFbdflkV57hY1r32K14Xvghl3G5T+OhamX36OHVyGH1WEBfmiOY5sxoG
23JZ/3z5H2YvAAT1hxflEMGnL0+yFvz3TlzmwfpBKNTTXSl/H7hH2q+nQdRA1LHY
Tirp0tthdiulNT/WbJxvKB5VXKYEmSrfBum5+ylNLQMEosyqrUbgKIeDJw7HZMH2
gMeYsmAx11jNcWrMDJbV3wQmbcwJucVw3kQ4QFoMrIU0trkxAOh/9deFpr67ldex
+GPoLHn9Xk6ZCYjG2wTzNZmkDq2V7oGaFhlxTnZ0GwORXFUxQ2PcEfFmEQzw1GnO
96ZTBexo1WtakBZ62G42iGD3WLzhX0BIClpC8YedH7Z0LQZdyB+gJ/GRyGACg9v7
iYBlt5zsl/a4rO3jhO9cJKjiM2jVLEvVOCHC03sbCXRUzzawGKCtreK7QCdJTxNp
LTAky1iRNNTELMsVY088j+5U0SBwEgrX5ZOOfMeldkHysHJz0s5x7X1kdS7ZgKZ7
AqD0WTKCV3vqBxQ+UZDWGHuAo3TN1Pt/obC/+483DDf+4vlVB6RCakh6A8hNlmfV
LUwctWzkd6d50IjA2e4hiMhURKZwpEjT4yTh4VIXfAM4jx1Ob6Dj6etdnOhv9jmK
l5BVIh8pZICh4VPl5jb1piIXCG2Ub6ISPGTAhkqYt/bPi/tvkfSo8SuciB85sJWw
h0itY+VDteVHTM+GwxqbMcz/1kF3YVm1RzSGGrBVsCrmUnjSagTc6iR4laDOBCzu
oQ/tN/W4kONi8tm2p1UaeLEfwKiIImIxasnjRgrFbN/siGGZ/Ed8aIoS3D3wChry
rc2hZTw6KeCWXPCJ232MHjnuHxuy3+vIdf4YNSjmI7w5UmFt/sLJ5HjAgkemeL59
Wx6cEnGvnip383LrIq2nAY7NQaATh/t2EYjAT/0CnX7XRljIJReb7Fq9Y9oAtuAS
Ix1OURoaWFW3Q4zIW1iPfT66iSiU/wYCtsto38QOe8HcXpmXxOoFFCdbZXlvKpm5
Li5+7NWoea7TRo1VInjogjYGf3JN0eRaZhrc91ezNrrhlIGrGaCogvdnAfRxtup/
+dOLf/CDRkvTHW4v/uF/fTSArH21+fooqHKRiPdn6E54eas4T1mA3Ten0tYG9WjQ
2m72sEDLfnYGo83h+zblR5+bXB3MNVMpKJVMXmzswmOKqvWRWvS8XIalrZnXPE63
09ys+qbPw4XTmLNbvxA3S9STXicEbO2+EqphyhqR7Lm8yqAKo1cy0y0GdOZhAtpm
cCBHer02ibR1ZPt/EQNnTqijlYytKPCkfrszrPhBG+PQ+ekx+XoTYlw60/0CbU28
P5YhfkepvzCX5R1bjM3w859kaZd/eTEZq3xBk6dpMp48Q8Ll4DonoOlcrgNnAqEX
Cn6xGqdS0QnjLd5nEJsIJvAVhx7XypY0W7jqFWdyiJ3xZdGcQadpfvFPtE40WcsJ
dD77Osoc8NNpOFXVFnU7FBhJ7qj6EPb02kJBb50ytKrs5saWG5/8z/pcq0DWZoTr
CyqX8aKBw79l9i0TYEwR4s0I4JqAlddnVevvzmnYwQz17pNQKKOhpOUtClMi8Lo9
2puR01Nd3xlEO5ZuPmJswhSzUEPHkIJ9hShBgnt7nCmnpgVrq5o9KJk8OmT6vAUf
O6mzhFJpCnUJC6IGTWz9zhY9AvIzti9cVaH+aRwSE3dAurhPfMQYYnCv7tZ9ihuB
AsFx5Yi8KjCcelbl6eyyIuu4Vn89DcxfyaGmVmATaZ06oNjxTv+wW0DqJPeXHPhF
9jtzljZ9NA9uT3dnLHUk1Ktf6jkQ7TFjtCUZvxysqEanGMXAzOSMO24m7ya9ErsI
dCxg76bW15Ff03/Im60KNYzvon/uPw/o8olFanOuDdiJUD7io211TgYTmM5jFZ6N
fgMnlc7/qui8sqStXzCozc5qbyWuWzIxoKHomf7lzFW/NIuD/7vPhBzJZjeE89i/
nnh/ACknRSwS6E3LerRHbZmGYhBNciTd4rV0Y/n7cpFKP/Kb0SG5cltx0JFV5MmT
J5NDUbSMcyiaOiTPMOpjmacN0cEjZMW+/VzYAQWdMtN62RAYAfoqopDK3jptEpGJ
+T710k4Ua4wGO4zm8QB5e3XLgkTGqYBO+Eza9yZsqsiQ4CDHwWbJ38j3zKxuijZy
h78awm1sumGRK+uGfwa6Yemj1hDbMgJgrvd8n6jzWNZKJNYV6W0FfmCbVTjmOMpE
kwtsE5jIqSs3FQBMlYg3rm07k0Tjk/4IcX0vAOCcLAXi3k7uKh06yttQjk7v22+z
g/nkowPXAdzrA0M9TliWs7GFoMFQDRYtI/J1Ffq0717zedv+7B6DMBYI3CcK1GkR
JYXKwyBcf4181Qtlt8zZIqdlzUXNrc7YeMFaeRQkNoQz708YBAEReG+irOXjuNPz
FzTMjp4RKnSdhdzvaML1Ynb0ero5zdKL/7GU7hSzC78NxqsOVrXNi0lfmYNn2YSx
8o3xdp7foFUKo6231CiHzZtzea6UVRlVHvp4Wr7JXlM42rPlzUqsYk54Dsk+YxaC
aSQuR6Gf7m3w2tp+0pWJ2VNGKHLSdS7Za6T+lCZ8endUjVnCdvsszLwqWzikbV9g
WcG29TjvfdZXiaO6EBj5MZhUSKyABT3VgtVDhWd6x1GevQFOG/gI1i9BSEw2+zIb
Qc43wKgl1MI3pvtigSyXWakVQBi2xFi03DG8mpDyO2ooSgE2Zt4vAbv9tVTanYBF
ZZ/cFi2VBZ30gWyUOpXJprF8LKAFvmsH9lCDCJnlDCpsrtW0SuzdNmDdBKcziZpd
G/VLHhzVJiVTcIyCjaqnfqNWSPIxhYqLCpqIszXj1iolVw93hxlCXDJpm5k0w+AH
j6ptClI0bt3HZh7Hcz2TtbFSU8bJu10Vmw9C2xfoJcd3022unuOxbFi1t7crFzZo
vl23CpFEkpO6QgxDRCA40LIgOzheM9d/kzALokn+nj88+TThL2LKtH/KNQyg7i7C
W6GY1q/F6yiQSF6aPme46CYanTe6sBJzjfqWsT9/jVNNWGSgcFa8rZ84G6YIsSJA
lzTJyt+XjWTjzvdazpa4DOcJrg6bjwIahFx8vScearyIf41dCW00DOLTYQ4Bscu1
oZLIqXIOslYEPDBwDrO8Mi4SwadzRWy6OQ3tyfp9ODWLGTbkzinD9W4ROukOch8E
vuqv0F+37qcsq40ceS6cSSzGUea7jJqksgC33U5pWyB5lHu3VijHZ/sTLi4z2W6O
aIC1NPGtlSE8vP5RBLIcLWXLlGVXPceVdJFzIopDoIZ/pImbyJ5GP06E3lxnKih1
RIHXda/PWSRwPUYFOU6X5RcNPcp5DTTpeqgTegdGYKnYDRxksdjDqhW/sUc81loC
OmfQ78Nc6ie4MUmQprNkdd3L/Qc0JCtXL5hhZROCnR8wqMfnpBFeLZ+CMf/BquMX
BueCfLR978u1/TRS8GVjRdBfTC4sMjQzT5jAJHIu9i56E95QrOTjBvvif/6HGRfe
iaXGPga2Y87yBXzG+HlZzLAs/eUZMYlGZ2fWGs5Un+0ARTOJ4UpMHJ/JFcOMSBdT
JiY06c1gH1bLdqox4ys/WT0tsSerk+yl3ZSEWYFosZLpXvz6uuOZ1O7JiSUT5yjA
UDjRXdxkBWf60I6XxFeRn2YR/UoRW9MmGBdyFaD4j7g+O2hVmZut2DAalmYGSh8I
W1udkr/YckltLV5s9gXfd6XcXbcIbZb6PX6Y+iWmuwRrm4uBnMqmJ+NTt1fsWleJ
pvWDPpH3Xws+sF38KyQ/H5ClWxlu/OSdLG75W2enH0Gs4oPVUNvtv87FofjjROl6
jyGMtbDexkCpscoXNR/TZCkqcW88x2/FV5nSdXJC7qpAiZ0tQ2ai0qYisJvbeLuD
kd/wDifaAq/ujPbRxAenP8J6+BcCaSp7cK6APRD1lVvBtPwg1Ct+kKMI6eAr0R6K
8kPRDQqkrZ0DbIxyeCW7INmUbqj0hoZcjPLLvJ/X8NDiNDGq62GHsp37GWLgmZzd
X8WFCJasyDp0ycCom3Fg/S2VUTBNiswW9jtp7j2GdXCiOIaaC/SlOKt5jSDI7cTn
lIUP6Wg34z/71TM9knCvMg9aOEggLLz+X2tBizIHKlyK+Vl8BOOmLsfLm1tlFM/K
0UsR3Om/U0rSgPLQe70YK1ix0zWK2Ovr7rVo8WRu7g1YgtgFdUhoQRWtfk3NyZHf
9mTOXJ60d9UBkDk7bqQQ/3wlhxIQlxz5yZFRDAXoVf4qnH+jJUm7JcGnMGUKuP/k
+Zj/80SlUPJIXX7RnBpzbTUNMBqOpdpCvejh3A+AkpCJdbkmLWm7VZReVP5UCQ9l
vgzXfhZFqLBNKgl0gTxDfqhTmd+S4VEUOsn4Rutza5mIatKSu1kCRKCJFPYsnnF/
DZ348BczzvTAKt812cKH77mjgG+GPbPB51QDzI0yDhhjc/EISaUFfFv5agUT9syS
m/9642iD79+h/RI/7Zva0NrZxRw2xLMjKeJPFGNuxt1ujIj5pfIuPfWdAqtNwuE/
X3jaKpCI2X6IS6ZTfUPC+iVSlBgWFQuJuFnWn1Ck+RoElmXdmHzhgg607qfWC5GL
JPmYiQXXl7pAG/QzffmUZSu8x4wW+FiiRcAU0AOBNkjUHYeNJrMtazJcAspPzBjx
VAo00S56naIG9fkXOr5OiXnVZwa2Zb/NzUCsLnthfnAGaz1yqZmiWARONNedsG0Z
OdrcSyW+Lka6qoEdAi+bK2CzNCMIDs8qpmawep4UWY8cZlOKjH6pKxNebi5APjlb
YLjAWdbR1/G6QNSP/3uhmguhOKu2teVADmZxaR/GMYZNtK6SE4+xf9tTkp2i0lUW
KqcHlWx0ygM8J8ezEWBkQRKCfj84rX6d22OwM3S+gPNzNzyRgHnEDP5WIAyGIs8S
csAj/Z1FKNM5VRCrfTKGYNQWt6fljEebqWxnj6eRIbHoYavbMrnRSoydAHaNS15F
j2B7nEtyw7gyzrnUVGJLZB1h9RO+7X7fHLoZesnaIMGgSzcUnwfDTZdl+vzmOcVU
5ZhvqEgi/edqwAWs0P1ZlOCWBMSzr8yqlw/VWcmKGo/MMBM6dKVWbYLycaL/1QKk
X4QuiQJgO3yWwO972hqI4LqPkOmb/6cQcrWDnk+itwm1hBye15/fsLlnZH4hYYjk
hEcBh8jqpGUQrf7G4VgNW/0R+ur71fHu7A+0mQj9OhLm09bxX3TynF4F4NQdxy0G
9hCnHz4JsNq+JvN8cWwGwjzAFNNaeoagvwYADTOJ0QFw5iWsavEorn6GXcfvOSba
9jsr7F9SU/2aWSelienGB8jYOYYvDTsqW7vzdrtcxsWcIvldtK4t6yZSoncXIgQ+
o+t0ZvPS33eH/keCM0uQ9nYWIOkuoVZcWhr/blZaySBtDrz473x/7LCWXivjvcHg
Tn1+r8lSfZTlYa2vdpR3xUXDNtmTNyk/Ho2q9Su8UIVAv7UR6KS6SauU195Y7Vil
wR9hoQOP4U/vN/pyT6iEfIhGeDmV3Z0Q4MOOWgF96QWB40LBH4eHjYZ+yeEqWmsX
aPkAD2h7v0EHJvR+VykHnAfllCypuiNV4WjcWZROvWlrO8Wyl8g0pjoNAStUUU2+
OGnCCKkXsQhaB1+Eaw0R9hTa6Nxtgn4P4yExqrERJYGRrje7NdcJpGVC4q2TCf+k
H6fmI3LNQH1GrkWvF3m/Tgpcr0xF5fe0DlfQS90cMcmLkh0WOXYWeay6hDpN69iR
1PDwc/sHPY1ldiDNT3LVT16lHvrJ3Q1BvHDguemuGlz6QG9FB8nFCx7kivrR0Q84
YUB9K3PcTKaGHLkp7FNJzOrI6wvO1Fmbv7/y8KfW10nKHH3ToPyQg5a8vviChi2T
W8z9uX0ZoofeWxDH8owwecFbT1UWY5tauSUSY+ZKs4O55lAivz9RTVKS5T5ewxdH
vspyrzEOEDCO3FWtZA3YnSPq3K5qBTp6dua2OfxqvddwpcGkrAz2REcjPbTblERZ
bxrsaQ+WrRqZ9N91x/yBtpSDKIwbLAb2h5iGGRtQxof5BR9lwvbNdr0mlPbBEs5A
Tilj59xxUKuE575djsKcZnFv5TriwR1V3vuuT1ku5CYjjOCQxv+A3pBwHkUTlVqG
ZDYvK7knseTxQTpkkBJj/YLoXdnCIUcQnWyXPAKCW6YXqgXJuY3/a3e8MWxNn0c1
Mei/jDtfFqlPLW0uLdDm9LI/FeUK7weujWqmE556WuDC0MCcWP9SGSD34HmR6ptc
E039gPrY5oqU5vUHnF0khvJxUTIZKyNgzAK76lO9B/EWDaJtXmJhEbewroEAA6UK
nNfv/gf5u6i+FPVGKhpTydWWEMnJrKtM1yrHe+6ubwMLrrZ5vcz8ZbaNyGi/DmnB
kUtug0phQmFfghUC8n+/kB4+Az0Jj5rk3RWVoGbd/YdpXe8wcErZlItWTIgeeHNX
MidFNwCh+nXmaWFBUZrMgUDiFfDoIgH3bpV0WYVqiLCkQhM4HZ5LwuAouMLyUYPD
yamGpEl8fcfliGZLWyu5cwPGeNnwvPzkmq4pgHzyCBQjIOtsMs5uz0R3wVMdBxlM
1wtptNbnefOtUQsJi3iRD0RSYl2wyhwyxr0V9eQqtOxiazyaD2hkxRtACvJcu+P5
6dYSr4fkf+YDW0ieKbVG+d7UP1VZePGqJkwyQ43YPQ3iSeV8vmxvkYqt+Ciqn6qA
FwaOjdFMD71+avvYwirUyiln5eMvGyJtXoZLfLUBTwcvLzPP5DOhzTVUL0xQ+uDe
ITpVy+e3gr2+tgZLZPr03FL+owex9trvcywHYp+TUDKb6RjWstpAcb4laIlps0KI
EOYjm8K38y6vBeXwullWUgkNIr+sEmsIKpyuO6cfAPGqJAoQ2k5w6luu/89iGxOP
72f0x1H46qwulW8kbjSRW0C/7lX08FgCX69AyLGi1FkldiXee0t+H4mpcrKPerdk
YbqMpEUnhIFeBI7FVcV7zDscCFvWu9AVfN5h9vrCVbhf+FmlH98VkEQI0PqTWmTo
RQ1VkJQINqXoeYqDILMRTJVyScq5nG4PztFCj8kzSh8Z7SHRhOqagjnGaidCzPq2
SOO+b7AJsCmuTfxISt/tEmd0ImnaR/pSp6F4kVJXWPID8yEPdIpL1ylR3QyySdzq
jcp+/K9kibVTgRA4rwftUgYh8SOjrJtiNEIqjNHU56fSRMLEvbEMKc2Vt3K8AHtn
3Ur0qAAITFQXDKzCM4SGr+Lw9vQKqLrcmg3jnB7EUN5qlatxrWFLI5QvC2pKWAgS
1+e2GcSDrKCONKLRoFfutRNW31cxrmGadc5eTs4gxaAfJ7DPJerRpflmz53s2PgB
II/qdTYaewtcl75745DT1bV7aySDW6TEzgPc+9/0ezevOGNcfYdQqFyaPPM2AdAc
lNVHiuS69ykYArSHrIuKjBZSIPB/YQlfhnU8HaWWfVhQOFfgmnmfebadlXQbKM7n
tStaKaGCpZdt4Y94a19poS4g/W6iUyspcGRaQ1xTG2jxzquf2ntqMPNjILI0QPDy
Y1mAn3Fku5XEpuqDFKfGvjXc5mV9aYcST2vowuK7d9DKXwHHhIOgNmchfvIDc8B0
uttwKEhCfDcTjbmqA0kvjsR6I+i8ipDPb64/PnrSYKCd05VRrGfzYwRWFiTz+l+c
eh3WjxAfsu1AQyhx4o1V/OAbA7O7CKp5ijYcxKf9sJs6FU7vrMB8vdyVV0XK1oAV
ntKUHE3DWLgzkYXwAdWkrmi4oZrRfPvYbKVLkPgQ1aPWUo6kRnR/KvdRb43qpKVU
6I6Ib3UfW9TKZPeWtERj8ioKvMhogsw0iIxKj5Z853D5ZPF9Y3nfgnzAEc0651f1
ELJR9/sq+wwxfqZ+yBcwBNG6I6+7JTVXFT3z7IOFd/E45P/67Fz9mVa/le82XU5/
RQVRPQdAji2LfPNjwQLWFMOeIGQEhpZTRviz4JIY3MBFRVBzvGa/pes0kwmCnDq4
5BkG+YwnMgbxOq3wGSnoax6+pu4CKKJxWCUFx9bw707KIkX1i8+PvqZwvlj2Yk0i
4bY0DlCM4x+9wIMIIllHwo+BljAT5JgCjHY/CZmJGageARtovRgQW7Wfn7GljeYM
NNSy+tLAKESzJArK5jgyxS1QXjj9/pqXmsDxFqf5xUaZ29nvuPh8PJTGF/qSPa94
Bs7cLzK6acjQNexUa2mOL8UAMNIElSXFiUuq2yZ6/H3ZFzPsMRGlIMVG7uo3bpcU
nthcLCsiSydbymGA67r/O2EQZpXICQshY6tyTBrbLu0yX3krIFtvGTd/z24TGmq5
KkZKUrx7d5NQu1o7avxgkbI+/sQoWzzRxLNke5oNTGPUDlUA2WkV7Ef8wXlCV0wK
KefXQYDVA2wNGXO+MKTzCD9Z9utQpmXzeiep6b8/97mJFcTn/ybBknle2iB8TL6j
X0EAPFKc+8ypN0haW1JJ9v6/24TFjorezynpHczXQoe56N/iBivyicjVyXYVsgqS
SBLufTxqlRLhXnR56eH+9sTReLoD0wPVCpZIJB005LBJdcMr7qAn/rmaK1WHV70D
Jqp1z5Od0eZ2v5ifff59ucHiMR0LZrS/h0F90iN4l/e00PgENtCqJgqZYhpsgPgU
r9K2O0AUvGWpwj/T1xM2UIkIL2MdlQqN1xYlvDG1ugZncV6mHwNlQdUC6icqMBF4
RSiLlPyJ/k4Biw6FieN2d99M+lZjDefFmWLtXXkaaGu7lJJYpVQXrA5Okd0FyhAw
fPeJK+JCxUBHcGR8lcabeXv0O2MZg7yiccfYCBCvehBj5Gykq9AtXd6AUdYFcvEi
sSvcBtK+GMpomkm4BnUtEQHrBAfjaSSOUdIFJQ2Af8xk0jNHkSNA1DjlHb3f0hXW
CqWJ6ZvgUf9P/1s9Zjb0mECs7FdI9e0GVA1gcNFLJyGeQjTFkw/AYtypkVMDn0ye
JzJcLZ1A4NsLr2iKqdavDEh5JskY1fqgitkaAn9M+3t9hOCnrFwiIdhVZ2Bu/LhX
RCLCZfWqU00NCHMAsne7S6kV+ct2Zn02Ie2NSkq4Ekcvz/+lqXl5y8L4Nwm++emX
Djql5eO4FfJu8/mwLYuHxyrhcabHfoCr6WljskhNIRWV4escjSB2AQX6gCUhJ+nE
DcRGiqK2kdCe4hcVfd/QpNiqiemPQDPP/H1p2tn6LP+PuFWUIa/edrifTWagUzOf
gohHBntADcU/32jG114zt0s4MvcPY6Vmz8ZPNnnDMIlZQD2xRJfdcfP1gXRaGOvq
tAP49RfayRBRu5EuIakb1IPDCt+Sj72irjN0pnu2X9GAqWp9GUsj9ynkP3UkU5ip
xbCm3PamIz6+OBFceYO3+wFAJpGQ46GRSPjdzjg5XdwOtZWjIHXdl+E7o+/Dmcqq
YKp21QH7UhTxAgiN4H9zv/DmnZ/rv4EEUvFbmj04oqzOtSrgcXkhu9zVZQbrACxz
twc9aanO3R/e+EQqbAonn7I49Kaz8WB9kb5zop8YOaSxdlpsStu728nd2V9FXcyV
3DiF/2fx0jyg4x1QB47Vru1MpiPWyWcRS+BlseZ7zQIu7yNnmabkkqC3UiSwkCDh
hoTa+XiohVlxrF/cOEXlpJ2vC+ugsfBIhvpqKyib2Kgx/5kjS445ODG8hajRQTGD
9WkLYP1pC78l4xRefahjfi1VAygYM6cwm2EqnAsGXH8TrFKPVQ285MgItKE7BISG
jhfMLoR3A6eDX7bJ0Sf14tU411FcmJUJZA/T0a49Slgtu2JVEcg8y9VmQEg8QqmS
BnBFPecZ45L+oeQcVG/w6/+hdlfcTn+4QDyG1xMoaW8vLB1NSuxcTilmByjLdWA6
eWiica5eKZSMblzDBgNWR7W+/hQ8lol05lMtv8JU/widoAYN8yiH9Hvwa85dI+/P
Z3+TRuS6vohWuTdgf48BJKV1FkD3cK0bS17LLdhQQahI2GcIgNsyFVXyVgV0sPKo
D3wzibSmIdtMoIMccKBtz1rCyYdtYFWmT54BNMrQz/OfjBtNvNZofqL3B6FBiwU6
AWptEid8XySmyyl4HkCbji+x35td7a4mvIdjKd2Cince1ghRh7RjrPOhoaONfNaE
00+VkirhXVFb+xs5akuJECzGaC38YO2PZQnP9JQ02dHDJtYuQBd8ybFGcYqwiOfb
1Vj0/tb7OWPUiYB7ijTiohdNNBoLKWpTQf7oiT7auOyd6r6z/6VKVJOaE/4LKMH4
QoDYZ2JjwGLWtO8zdXnuIRdOKRNYC25pJ8NpNZIcDCwWbklUpx9inNR2idfovB24
88U6j7531S201k+rf4GD3t3dwxJN37EDNO4mB4fDdsviW6/sLfRDGQkGA+CIKJe6
2/OcZ/EUkiqjOeuzCbCiv4YyuRrqXDn6+XLq64EqPwyztOcx67/sHisWHDziBEIo
1sztLdFjcmkFhuQlc2yBGSGf4BZEvAWdS4rI6U6obgNVf3nSGz8deIPf8f6680a1
o9xZCDxOagYat+eT7z+nfswdB6h1Vwp8n8B2JiX/CSmSCOdVnU7qgBjNHf1h6U2G
d/P5/Ho8Sdr/CoBU5jSx7f2B8S1j2Z4EgsIDtAPHFzvMLQdAdXRhQKtULpZtS5vS
2AZCUPAfxAzpf7sT/LJr1GqJsiozcl4vf95aTNLBdd/dEHzblW33UTLd7E6u/iTz
2yr4lfeHUi/eCgsYhz3OHV5W+5aP87fx/8qOI8UdVS5Cdpbbr8mREByjjiRVl4N1
3NrUQoXgLOgAuwRho386rN2Sa63j3qbNUPYF1cFVMHRYr4Z9IQ802XR2Kn5iDvJe
ofb7VuW3RhNdlxqK0XWNKTVvqZFEllvkoyWzbn8MNHz7lhjHMD60edzv3oBLWYzF
BnpXRjbq/dzEpmbS/XFUOd6dB3wRTeJcVpizWmrBoWr2Kv1+ZEBcRzZM5twNyn79
rlYSwML81LW03hRcGywrC73mC0klPfAmFy0/vu7auDAP3SmOwoqjcQJ4DeA2464F
f9zbLCKXrR1edGx5glpEy9cY5poOiM9smVaRZAifswyPPDZ/CPH/a+VWLoY/x5cJ
EcARnPdvC6xZ9vDLm2GXfu/wYgrPJaBnlQYz/VLDuW9hJ4qqRBmOldflct4u/gZm
AJlc4dpr2hbL27SyiZXB4MhehDzgux/HkC015K6Bw6d15zaE8NrqN0wFEXMRzmRx
e4MwomjuCjyaMwu38ty7621r+tPYlxJ2Jiv5YPYUNuezHYb03zlrsy9S69SVTHfQ
znEA8K2cToPd7CcfLd+ZHoK83bMlpj8E2fcpgQ9CxNldf6bAeKvHz04vla9sJWqO
5M6Nnr+jwlvvYEZEWq3KnXUKXJM/8ye8938hj5HrXYQQLvQc9xtcm2OT8numT1Iz
Oy0hXy1OQ/Wgi9NdxNQvmti54EdF3KEhNOxbBjbHbYtJVMZmB6FuTNGysgc0YX/g
eendRqRcjIXU0CI7wi8FmuivKLx+xRS/9FTv93RCNiadpZ9C9Yh5Y/nwpOhpUVyl
x41u0NeQWUj+ZR1wKDirlj4//Bi98Mll9iH0L+zj8e3OwESx3f38AO1/RRYWAC0j
AE4cgDWME0awbSAzDQYu3Xc5fj5cEwawkgnY2EOlurU1O4uDt+BZWnbMwEYPVwSk
Hlj5SqYxO4A5Vy8yNCTe/+ffShATaGtSYo5+wxHjG2aDU1/UtMKHswPM3KKuw7Rq
8kP9ghw7ZG2KTS8aAzZMBtNl+B2YUxK/w4st7BjXWo3+3rMJmZFj85BNpiq2XFJ0
HtqbTXr6cdAXHjZhy769pTBJ9sDZ91w560XFV6fdTJlEld7/xuRsqouIA+DdmIJa
ERT3VBEb7AS5dscoT7Nv5srZUbqvx96CRC1QBK5tLPfNPSR33/VmegC5VxUNnp3+
0w/qXoQou6IxU3DqlKSYwq1iuXvopAl/Vy5rsQWMK6t0XEuCW6X1z9iN/U2Mfdkj
XhlHD6d06t82egKe2bDN2sGzs5tC2F8fRg4jbIJbHH66ssTF9lfeLGZI/qJcOW4J
xMydboRib4lIINYl7iXrJFwNMgnxlZZbjSiqPaue1nNKwAXQjwZU3hu72vx04tK0
959cEADj0PL0wuhi64fe6n5itwupEfZ1dv6KZ36JMILs1MVRs2CVfwiyfrNL6Hyt
6alqD4Wr8GFEyp9bQoD8fdYCugoQmqFY2XVpWi7uEmWcL2FdDjOPK4RJYHzsbqoj
Xs8+K0BR3PGRjISRKm2xa9zF3i/J+Ac4jhYUUNVya/0nzYjaN+X6sfcQBXUwnU40
gwx7lrBE1O/YzZKijekdSgHn6hBy5Kn8+0dmRspSpp+5ZY7tVAH2FwysepIecgQr
eUaKv9j6IqG9fkGpMz5JYDXPWmQB1McDbDsy4+f7DyjV4pIy9NopyvNMzardSon6
iuikm8Lf1/zBq3yoz+kuLNu/4LO+lQerOtH6Alakp34b+xuposIql8ifazmsS5j7
e/yRwLXR564R8lXgA8mmZafnPyVnD5PFWNYMebEwVJtxdIcEpd7PKqEkYH7OGDx1
y2MD+xdc+oVITotT5/mWIyU8W8zjoeLQ5mYWL29jZHcJ4LotWwT9lGrlGNWe0RYe
s6fgHZdm6cXnhf7WQz86O3euXNy8j0da+jujBtrd7zraKUdf+kYNW5RXoV5wol2I
4sXXmRE36oYerrSrOhNXNcVuRA8oqpqxPS4DMRAksAOQpa7WyK6pzdbX7YBfDvXm
OCCmyfEhzafRP+Gy785+Z9CkE5fUOi3btDDjkRQUDcPFJtj4F7diQSJ/z9bavl7+
mWYJDbfMBa06SNEx8PElpsP4UiDLjZkQRjmahW1pQiZtIb75yapRTUq1fjTGBPcs
1vJOnqIHEgFjGACxBr38zQenuf+UKRuKF7pYcx12Uzjjmbz4LX+hHGfhZSqIhuTe
7n6LXgWFYhun4WBIWixMygZ19tWY8o8ExZFZcQwFw51gp/yP5dVFRmaMjGHxuNCf
551e1ua/H4hKuzFh/MpnhltmhmwOK7yJJEmAjW16ahpM7GJDw7O03LvpzTxxIp/s
sy8xOaHNe+BbU7sJCYZruQ78nghhuu76HsiZKQMI5n9r58QnaQcBzujZl08TPwQm
uv2EJhiwRx717jTJ3ivjFQCBubvrmV7FYiwvKvwOADqibNcYbppddD4Ar9veluvg
QUpFKlhDoSHlcmmqoxQHYJR4ZhS7IwpdJIAoyAf1yyer97j7zKPm3z1FwrBFPV4O
AfqDI8GIc2xjwzh4jGXbt5SaaX01ax7pt0uAV5P/sssBRS87rMoJ02e2qgh1TrmL
dtwX/TZEFaW2MIOKYIsz9vEx04/qkhUsj+MwBtOat9H5zZCuqnoZyQ6PLy393EJN
39q1tblpp/S/iGi/rInRxHdDyr0A4UoMYdKIQW//tRmiTGy2GRoswe2PJuf8uB4f
LzmnjsR+yTftPSCw7CyWw07/2XauBLvjauQBX/roiN+Gkpc2KyRlSbQnUxEpNNkj
+mtgYnqmy3f6ERqc6/acoQ+ujQ77aTizg+Vnb/hrhDFIhyoGFjkq5/cfR0nQ4pxs
whMqgY8v3AbFf1seVQIG6YaIa46Cr7MqA2SNZA93PGNCMV3Er81U2b+NWhAoa6sn
9nTu0TCupy7vOBUPzT7XpJmeITJZzsFnclCcyLtBuC7WViNH+0kECJqNrGDVF+Nt
w2ciVTdkEaBjJ9JJXvVY/ujPSDZuWR3E0KvKZCBeFOOzlxTjhmGKIflI2Lb90MLV
3si65t6PU9UkLKgsfnUAlj3OoJLR7AR0j9I3gl4gmxyzU2Y5hlA1X1foC2PNTlMS
54Tgz0DrxIXv6uMZTHC/uwgICz/ILhxubs/fs4ovO53TuDVgHDXIC75aZ8DrbFIS
disPns9PcPJxCfANobeYAVz6eyTxluJIfPRLal5mjP+hFRIDOCwqckQeTe4X0v/H
e7Ej9KjtvszOR1b1pYR/rBaTEpS/u1mnlXEvdGUCZx2/YT/dOXdTd74+/j7hONbC
U/4qX/9j7DhxfUQYs6a2zgzva/pVQSydeAW20Rn7bJPkBkmdowHnkUGIOdGbpSNH
USIH32ESuWkyU/1+V59C/2QhYq9LrbnvMPhKpeHciQiAOyY4EgPz9DDh1c4Y9VPq
YGDP9S97Yyr8BcYEE+doZ6PS+K/jt4fJ5kk03hX6zQEAGz9TiYpdwBcqNwv0QNkp
KdNliYMbk+qVbzYaCCDNZVb0SMo1SicTYU7SL9/+z0r7zhhDX0+02OhAY/8LdNNs
XK3RK0zhUpEnPOLiG5GghWeotWWwNQt3VjQORa8/zK5kMsSMhhgyevw9EqZw98Q4
bVsFPXdYY6OOZ4xVf4hz8putLSrUS7GGj0xI59g3l+q3vEJqXSJcP24GNI5k7YJF
RVXn6R+30Verx9IZ2WFlDfkXRQFPOWzbLqgstQpDssnRqNNy5+69SNZO8yRo185Y
09Zy8WkS7009fjl/vdkEvJvv8sf0GsodgLHkea/g4FHYs3O+I1Xu+c0iszYJKlSi
KYj8KBGdWeIRueG9Ok1GZiN5f8wHPFS/ehw2A5GTLP3e7uFLzkVeODGQNC1li7QL
WSvw6H4gGwEQqyrp8byq1R8XlYHMKlqk+srmztINLS/P2Z8z8vSuHK4dS0zeh4fZ
eEhrAMU2NzpCkKFkr/0yEZ2c+SQ8jhsedwFCA8+XwVNvOTTYrFssbWDu7A7mETna
vb9W1kKWtldsq26kBQkK3mqzO0R9X4n5sy3bZ/rw1ituzZiRJjpZ+deYPYBnINZZ
285ycFp/kT015MK+ufY1UjPD3fv1Pm2ofWIHQ6tYIGILsDW3mMesCtLz5xQwa1m6
/tA5WOC7M53D56UETprDr/3F75R2OvezFutz0MZT2Gb6SzTXoeDJJxpD74P9858u
KtcVxvR2WTK9jCNkCW2VqRW7mRDIf88typleqFhibv3x5VQkUoqLfiF8VaHHm4GU
DP599eNjmAfCar/9/eSKd3wtTtctIdPHp8KQ29hV/d/LT1Dq44Pzw/UOfg8/bTSS
kz43/VlrQToP3dG2QSL/1rh1Hr0GtrSsBTdkJ+uPrmJEfBa47XpnbBSBSWQii0KZ
aGgjWGBWdWnCuQBD5It4TYWVHwpy875wO/E1zNoqmVdyRTCwe9P7PxC2YG32c7ge
VPavr7kLhYuxlredvOef4R3EmvgpxYMHbEN6dUNBAJ1aAupsI10iNrHbHZoODouM
553LWspKsAfo9hJ3M2Lnblg257XSM9u2trhcJkpugBzvAjXLG2Vl96gRLvFdNkh5
k7nki4fXWGTVbrYUkpvjOH9YjMr/C5N3WIxNW8PeEq+vlEljzlkYC94lYejtwIWk
27yJ8lN+NktMcPg8xQ8Ogyq/29yPHPIvo8XcrT6z1kMfvnR3IgfATf/bd/jDRuyv
XYcOM1RIsOOyALraJq6hX2q6UC2ZupC0JinBu52eb5sW+yyFoHH0HJwqPS/s6CN1
/w13/zRzyURnYTntd5J2sD6grV1BhRpFmYRKTcbmsOCQCgRn20ULhMb0WEjcPO/1
r+CUa2CfeE6aU9WEyMNWNjyLiI7w1S6STfIltqJFxbfWr/1zZ+s2dGOJN63RhO9a
QF567hqz5pdpw1/6fzxeUqVw2Skldloy9nemtIenqUisZffr2wVNFuo5Q9wNpM82
2nWf8DJJPf3RSUf2+xwJGBGqosAgfIxdz584XizRFlgs3XKySJHHoo+0ykTez0HN
igdGvweDQTMKc8xnHJsnwH9NU1Wiw54csQKSd/ScTJECrcZcnojWyrAH9X9PEZYE
SzwVsMBBZ0uNVHZnniKFynJaRyrMuvLthUFxyPRO5pF2sgaUt9IWQQ321SM3rhnF
FEiC5UvVButcI5y4i6SFgaYLNFzW9xmBd5WC2MWqY+0oCK/yIoVk/k5q/HKoLnmT
66frUiptyVU1SwvhVyltdFE2b/nlCMet3jJVhckHPUbx5gqVkDBEK7h0v5IU5UUN
T5q7/wEXCKA1ucP93p4K0QN8UW26k17tCDHkna0usZGD18MSXy7bt/NM9Dj7XdfM
xJre5AIHQTIWbiyFj+3AdUhVtpDeVbZjZ4uwMeyt4vcU3x9ii8dzTN9dy30U5NV0
zwirPFcuz1QKWDE1tl+RmCaZUVqDL606yfgVL1yL8T3vnXr0DtOo6hYj/8CyRq/D
jeZ1G+QBk8wmHSE9NwNx/Qc8+q4Vo8ZkJUxNA7H1pDS/pSe+balcpl1hCZIMQ919
ecOI0uDVcNtwyhc/UpUGLJUfMusVtq7qyPWKlgQj6/WNH3sKwC9nzMleGFDf4Ntn
3tg3SUEuGtLT71RRb6Hk9Il7G5PT6zCtZGUCUIXKpdReujlWLtEtG3PC6+b6dfS/
4Xp88KtWdVG69W3r1g8M7VDTKIvQulnVReaNSrSywdAhNWIvTxx/eq/i1GnLE2YL
tzcQcs/cZR6OgZtzGq36WbZiI2woR7Zp65HPP+TyYmabhiHuiiqwv47LkZc6NAwR
x08YgiyHvrRHwxKqn9i9/UCNJfVrBGcsX0x4GAQkNwjFOGxfFFMmMKR/jBXkfQ98
7KCYJBCIkCeLD/+ptf2PxFs7NCWCn1MdImbGtgrHrQiekdIjWRsV7kzrrMYInpgG
TCkJYnS9ezbbV7jd7iVVjKlSiGqzs41Xhauf5brVK8W8q1xBZ0CrNDM/9RON4yQx
jGc/8/ybB3BdKtJoSOqTwU1ebWWJs5D+SNRNYNgpCim72QyhIscVaVmZ+fRBp/pT
EEV+3snRVAxm5wGIGHpNOQeMYKsKGcbrDQIOGiZlKff7c+XIejS9gXU5QAseRCHa
UgqS6Pwubto6CF//MX5T6C8IWVSyCihcL7qME/Wjx95qgl/uBgSkRb5M+gopCF4g
oarot6KkPrOl5iz63alzUtqbYty3n8WT/Ik/o/lohDxJO3NsdJNaQjPY8i4uWoEF
mqFPEBXytOqu3FfvTx3NzXnqkHVRo0H7JrIBF7MkkF1hdH+7NtZqP9wM3w4vfFGl
2hGCgugfBSNMwwSLb07zeU23MTKi5nmKhGzgEI9yL307g6p1yIJqtevXgBnr2Bu2
ZLCJ5aDY+bPdVf+MX5JMlJ+/WCLAaJJRL/qdMb/1jIbsTc+GLQwJaY9djJXETR1s
vViANQ3cAKgQ4yesznphr8kdOBRRVpor5aQIdNCz/y7XPt9phSKkRUgJRpYqWK28
8AdwhyPmh72wJEnis9NJggdXkGoyq/qWoNNZgaLYAlt+8CTUXVRsQww6MnfbHcaq
3hPp/FafmGgYpIGuy9VV+CdEeWrvFOgdMgrWRWh/udIjOeSeJYw605+tLCpWJ60X
bcYjEMVHPDXTDxbkKe/PMNst9liWRbKj2CFlu1uNZvZiM98dMwlv76QsYBDxGiMD
OBRD6kbetN+pU03jN28q7B8Bt5RPLt13gSzKpPgLOW1kg2ttFqU/g7O6n9YW0F9F
xf7EkwOWitVqg2iNadavl3SnHUPsHF5SjMz616IIXYFs5Ct2ePInMAkaOjyVRTL6
dTB+dQU85xB3IQwOsM8V7j/kkQsT+GLhVaHxPLilPphYiSJvFzd8EBEGPRpJYwqy
zRjtKGmQXe4Zlj1NdUhN6ebi/+qmhpwFVHJyhkRtYIvNEul3AtgolO5wIhUdkd6P
A/bPs6UjrOTcFJ5gf/LvPXEQ8t55mS7V6Tb8VCqeF3dIqKNDaEy7+ivqIVKa7L0d
tiHt96WI9i6WgBN40x+oK+iLYqeQHyUMjCZCDAQgqnnOWlLQ41l9VPXmc3Jmus0v
WZVH+ELE4mB6kdWT0FAlSJpBpmkZq/ZqR7u5HFPwBmZLKK4ORfNb8PO/IpljPnnK
aP8RxaHlxYu0sDUefwu4VY2fHZ5o8Xhy0M/tFY5kwJTArO/dxag9Y/bZvPbBwHIn
icrMTgP4vBGvsvZ5v/EBp8lkmT4Iv91Smc4T4zWBvMz9yc+6pPkg5F6nsfonem4Q
5E7E8ha2gIE0uKDHyd7m+Lk5fGyplLGxyjz+qczGR6gQ0MoX8BFaelvRpIVncUeL
8SDfCSLXQ+NkwtiTO9sWuyV3kCgVdyXGNQEZYzXAyyzPdavuxOH2aj2W1kReDiK2
RNf3XBUnEFqgXcfgt+iT4MwgGpyWPpW4lb0mVAzVhhjrcbfx+8dZgKINQrZqhhlB
AesNz3VFL2Zg4mzAaxuNM1Mf0mo6kfJESirJe2OkRjkT4kFTieJj8TZFgAiWi4JL
U7HuWSmpGRnzMNPVWNhv1aPvRPnfINAEKjiEXWj+DL7JmqOye6OXodoxpw8bJ3u8
gM+VAGTfsNop/9on6GFkx5phR8yXYm2xA+ViwzoUWuRuLSlUC56YN+5iploYHFTb
SL6a4gSkkNzBQ/E0rhBxE5gRSgmqN8T2lFneIUp3x2Txr/IbQCdtn5Wf7v+u1lUN
Ct7LLwXZT9XOBvpsafDb8l/VEnBUD4V9w6cSt3621iIG8q2sIesOZ1mgNVpmG8XQ
BlcBUu593OsafeferFpBYTm/M7fbc4OJ+/1XsdAUCNNbbtbET+kGH6pQHO1OpLfA
AoMnjPfmEr0BKECQcSHRxjBwThAw/6ozMPuXPQfR+Ug2u5jm5iEezow2PAkdGEAE
tDN57BHIH0L8h1qrISUJcJfX3BfOpnpl50Lnf8SrVAOpmCL2N1YzWbbzo1JIt4AR
xeTJv1a830EFMkxdfRQQFP1IbynBvH5TIVZ9yfwKfcWJgApepxlTSYUedU1C/06j
HFKq9mllpg2Dabvzuwk2APPUQIqlBPuBjaRj+WpGAma+yV8J+jWOOqU59Sc7Gq1x
BeZKfAUWV9s4MYF/blAmCZX1Tn1/TlZCwWepyF+h/JjL2xFEre3orVEa+BSmmd9B
ytnYbXwOPjSOGStqhdzogq4iC+YtWrs5mR6+G/GJH1238Cpb0WoNnqPht1iwbG+Z
lnwpLSL4P4ihtSGp5ocw241Vslz6t9NCHFHG/3AN6QbqGs4/pKpklQt6gOp7KrAt
FgMw8oOpXazejfo3VpH+em8MTpriZEnji/+bvtFIAbIbK3g6wDdCUQw+vU7v9J2k
EaxWdSXTK3PdVxl7D5jdm+E2jdXQoGMQ0b9vbHwPJAAkQGxlM+cYdvrt0dC+uQrs
5fCTgAmwvbtXkveDN/ggX7d2Wp0bdHa1bilGHnxcJ5CZs4awATHbbuW3tEj3iJ4i
Jh8UTKSoz9nvswhFvFiQwkh9W8TxC2pk7H5tsngeTV7XbbZmhhwrEvSBiSxSW89S
hlNceNpDlLvqR/woeMxnwc+Lqw5JQD1n2fXOizBVX/G710SeazNK2GwzFyKOgIdz
100tNmzuCUewZxcGHeb1RyF1wj8/OqQzBrxh+p0T8NRYiGQyhL9QpW3ZAZDtXf39
Uq/CgH2g7WHlgvPm/oKlnkkv9IwSpG1elG9tdZtB6jRrLQFxH5GGbW+4KFtyC1P7
CJ3Q7DvXm/V8N3Qvux2ZDG82B9KTXpX9JemtXN/tCON7c19iKu9lJVSprIblEcMn
0RHblcJTmml0mM5izwptDD1NolbkKNhJIvEM59MFingh0UkKjhxlir0FPWjhAd5y
FNXq+C0zyDMDyW86MbbNP3YM6dyIbWbR2Wg9IvehDzfFnsD3gN8nTGuTndEgBa2X
+F1tFwY6/0ZhWL/b4oU32sBwyk0aegysajbBl4yv8wrcr4MWICGllQ/3p49dK78i
TuXgutzkYX8uHpulorXfVjttjoMWKWH+u3j5Oif0sW9KWHX48auhmE+4MZBvwFiw
cpfGvKuN6WPYwwOicrvLdJ/q3HPksk1W/svdb7/2mQDS8gizBHR//MCZXqrQj+Hm
nAGp2iC9axsWXQ1NeUFb/5h6B8FeiFgHGGCAB8or4XMmjhF2QhKXJAyewS3934+f
RFKZ71pICJbJ0A7Fpj/KRyB4Gkt1bMLicjJ4xTCZm5tFZeit5h4kLD049eq9kav3
2sFUWzCINf1wNR3rCi5VXyX/D9DYMFUQLZ6i4D0UisDc5d/soIUfC3mgdJIqyZbJ
SGaGLGtyThcXGMKeJhobNH8j62x0PLs1LIrB6dlQnOM1HGJ147iuyZVAjdh4smPz
dsFG1yUCIOxPa1jCl8HA8JOQTxLxRoQVixASbMdgj4WQ4gbjo6uCcJh//7ThRx4N
qz33gAMMYmOc53ADVNq4llsSIbQJzIkaQZo/Uc6M7CjRMZ04a0qQAhDGBzouFqPb
ar7jGz6zGxxq4T7+TPk847G4688oYeF+Ct0qOdMlkilFYoYuxORmO6jWAH5HeoB6
x3dtmfgGi7UfWiwK8QjDU3m+ZFbD9bRONI9cTn1/2szunQq7r2O2TsCwB0lD2Vx8
A94NEvQ1LshtrkPWMIC2Z31GVV2JUXpmdN1ddw1SXz0=
`pragma protect end_protected

`endif // `ifndef _VF_AXI_MSTR_HNDLR_SV_


