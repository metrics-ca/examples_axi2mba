//----------------------------------------------------------------------
/**
 * @file vsl_msbe.sv
 * @brief Defines VSL Memory Scoreboard Entry class.
 *
 * This file contains the following VSL memory scoreboard entry related
 * classes.
 * - VSL scoreboard entry class
 * - VSL scoreboard entry map(associative array) class
 */
/*
 * Copyright (C) 2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_MSBE_SV_
`define _VSL_MSBE_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
oQRA8egg2cMYPhv09zN7Epl+xN6YtqG1qXgrDkP7a6BobZNBv+DAMNLufnfcoOsH
TKbbyTiT8Lbyz1oKRpcOsDuINHwJE+lz8N5s1Zgh1S7NxqLthQe8lmOnkC/D/Ejl
ZSVhEVHWtPTu+mJXBOlsngwKptT8Vp2gBusb2CmGZ7s6dI5c7myUN9NbLgPSL6sv
lP3zjpxsUZykI2J23hRWnDgRVPa/NjPu2dZ5mSsY6estqo3SAcrjS4o6YadyKvCJ
vP350pZbSTRQLIVhl5u8pUA3fc84avb6G2PjiUi8xNuicVVG+LkpXsKID8RVOISf
rW98jX7qZuSoG11x1uv2cA==
`pragma protect data_block
CNRrDQRf11BqmFADLPyBsGvx75eINE6fPJT507Ep1krl9TLF/+GkLSHEfUzf/Ftm
IwDDn5KsSKFG3IzuON0eGSbYPJsFJHlKTTh0CS5aLpZcL4Tc9Hm5/DqDdCDX2nRW
AZaVKH01RKCDJIS7M/Q8ISYzzQyUJThHUZlbEURrM+8ivMVwxSubeKfeP6kknMLe
/tUQ63NJDPyJrAV5D4Gtmam3JOLGw/LYe2Zbgp8apxhK9Q/AapVTWhsg5UanlFhx
NrZx6VjLSgCSbnH6xfSY1YPMCvf+NGvpe0ZN6qQzVDKl7POTVPZy3sOFtaLGIUW9
3iN+dSYRAh+ibrHmYuOxgNh7NC+U889uAKmuOE4+i27RxgIwY8rRYGe0OGlRIvyy
KjpsoRpme7IrvGHk2eCHSEHffhXXFhry8ryVLUwVeJs1vgioiJ2eGFnTSoLTpesL
7o9JNmZpCfZUUtblO8I5m5qWF4VCjIx//TmiXwpDuFhKGPijjDcL0c6mf7c0hSSv
TeL23yNs5Tum01icjwvAqXIYa/jp5gwapTeUSkoljBzO8uom8CFOjwlTOlTTbBvD
lFBvBEol4O1wKaqsB51a6H7hR8EAytJkfAnYRVOgPoREaVzNMcNgKaUswQI9KLCa
Yj6AghW2a2hVbXS7KV+Gp2T+9x8BYk1YIZn1NlbnX1ixv7EyDe5ft1bHrLkyKP04
JnXtFspdVb36sqHUS6k+nDscf+quO1exKvBwZ1WdNJgqKWRcAaYd6jfYJgkDudPe
z6m39BKQItnlCsbRVbVgpSa8eooYT9wBY9s9QBQr4LIu8jUj+WK9CuhqzpllkIYV
NcQUqMkSP67cSx03FmUkCDKu7BzF59rZiLlBQnDStRVoa/Xix3Y+YjtE+CY4wO5l
FkQwhcuec5NPQz4L8sKsV1PW/EsAbX+S6+Sq0elc5GfpdranCsyHgLVxl2m/xCf1
aXcxS6Azvjbxp3KdJJtfvxB1ZpSpBjv1XZeftsZ7PceSz8whxRv4isiIlvte2K1z
YdEYhqUSJqEAsXnPU7Kruna/e8NsRIrCODU8Ng81uCXHhYK8l1W6xoRGWmHQ/KTJ
WgEy7rkzOJAIGbOSOQ1cCUEed5SC1F/M5/IW5wZF6sUHNTl2MqnZh8coUJNl3KbL
Cy8watSofgZHOgADsZe15vpQISZK+yEM9EfiWb4SL0pcSUv5fzTrg5HksfeQYO9/
MuWi3E2o57eZuh8q4j383s6T8J2V9KksVwyebbB8SxPQEKA/l4Q8kkR28iC6Q8gC
1FFngsCmPkndN5ubZBRiji9KsE5Y829PuOx0iwizlLqnxHj69Lu6m2yP89cEiBsL
ouehn7d55U4RwHg/F72hy2LHGaIGzLuUx0S26Y44lqqAF4hV2UMwcmy0w0YJH1NT
9n7fdIZg4vkoOAR18EcDsNQyWAK+x1/h1TacU8arYUhUFlMjSfp3wFbEYsapK7r2
NrlBoo8h1c4SSxdcWK6/8tZGVQidlx8P/xndWpN7u5NdMRHi62nAjOo6bWgJaUyn
X3Kep3YfCYS0LVvtVZwQBYtJVF552xl7T3lbI6UHe5GqdJ8uPR/b9awF6lq39nMD
vzGkJnuo0IR2evDsMlQBlHWu5nl9ysjVB+6vJ80938hUdcjX3ZFh+fCMAVsgup0a
2ftmsMArPhnyCpQTHR6a2uoNZPQ3yHKtbkZCCvYhZSMzZ348wNBUJqdXStKyDyJi
rKzzLIK7jG5haNtVI7Lq1RFP/uNlp9AFixnAWeWMgP0DKlUPmAXLNIUIWh52zcEP
BUG0dZ7cRMeWYxwtBa3i38YpLsrMDMLVl6f5EPpLdbTpngfLgKtP4PjSMu+Ww0tw
a3u19GOx1SHQvbZgCOCvA+HQBRM7JP4/1zBxWDv5gcqvkkIwb1zPPHPjFh4fjfxO
T1U/27FHfY9IyvGrCDBOi7n8ZueJMt7IUF13iULr6KliyyH0FKeEjJqL0bA3Du/I
5nu/T9R5kipcTzeiLm6phZVe2qAtKVjQvAJChKjxJ5G/hNDk+n5tt4nDFhjASC6B
iX56pt+pRoFATANOLy+GdGOFgeVgmJQtGbPfW9AuHjW5QCFjnZmgFe2k3gSraeLV
UZFfTj7j76eepaS7selqvWX79I5E0ZJo2LyHrzDxgs8K19wR2h/nunTmzBkEcMQQ
5TxCbkdy+zq38F+qbo2h77AFpIiWy7TQk2/jd70bWlQ9Ecd7e9S7/5w7lrZLUcvI
AQrLgx5ypdDxl/1MzWejHGMNDinIQHdeUU1paiXQgfrnUbnz/lLjJrwSM+JEUItN
CQaDVQdooGFY59hgwHtaeZLqVQlXCrKjtozvKGG86lGF1eUC3JM1+vOBoXOXI5uY
wQbT8f7CEBnsZODPC5WZTTOp4rEWxEtKlK+tvNo1T+xFeRjiq+od2lpz05yueORt
kGWDAHZq2nANykXKoC7AKIxnFEpgX5pMfzTH9nCtjqgofZvcbruBovmSwmXxQD7f
uWvVZHjOMRLp2xEyU7MvpFpGljFnXumaukbrofngFivlSelf/wuhcqZ9ca+d91rj
967xPN7Mx6asJVsxOjWI32HSyFfaEzeJ4a5WSQZU8Y3xxY5n6ye9eIyi3Zv+0uEP
PuqVhkFwtLb4wdjucZauv3LeOGBgn1Bp7uwtg5R+wyCtv1DcTw4xEu5EttoDyzt6
UWCYXoj8Xtz5ryQWk6kbir8jvhm3ET2koX8oeiA5t220JSXTWd6qzlqR8z+8s4q0
JMMfieXLx+fvlfzKgNBnKm2SCVnT6K1pyoDGe8KSWTbpPf/bk9G388nOxFIYLJ1k
Yq0kPQuXdpXf8ZPgzoeJzOLLAktWb8FADys0peAFcVJUGRdjPBc+8Xwlf4J/0e1U
n+n7el3m6i3da0K/f5YufHQI06Aqk+rHyiJzTaEuEBT9sptF628dI1jSfDXzykXt
Ja1Knmf8lOBFa+f6/z2etbzomu7QoE4Cf1W6TsRA0NwEddfYTPoprRdOn6CbK9wR
FT7HL7YoXoN9Dmy+JueOG/2uuVJF64gCzgNSu+HVOe9wtvSQKlJvbL1MkD35fIBx
a0qSXheswEo6pdAG3D7N/iL5I3k5cMVS8FM46kvjfdvu5qONL3gWShVFyXCQWEP/
qH+MdNMRYkzi5y2X5LlGUgdwXNVu+ukUwVeUI46+D3vFpVniVDl/DtZUjXhqpGG9
KnxQPVDBkSOHDUzoPXm25o0bKNoNuHuzhuI4r9CkBXQQiVIcSV/oJ00+aYEwnoHv
VLZIKmPDPAtKOzek6aZGIEPa5gspnYtoF7KDj0ITMRoNJn5qg8Kt/thGm3hytlbp
vTpq9NhFMj543zh2RytQRqj6OswrWAMnAiWIw8ax2g6b1NJfApCtzLFXqE0nBd+d
gebYWi7Mpeyg/6DAhRDRM747ashSph68CJk/1cRkh0jytJCmlq5kdtFrhgVbAnkk
CG9e3NsRI5CrVnXB6VJQLNioEzNFT42nHWBL+2HUZKzgs8XZlW2z6g3QLV2ezMZL
vbgSI+0yQFzA55mn3zXoUcmWFc8FfNP1JPGhP/tXietFWvwdxr3FssQphjiJJv4i
XTxVJaIRM07KNpQjgXMA5vXNgCXDmbBFQ44rj4HM1gZPdDwIgcxYQTFAzq5m/7m5
Kq6BgbMOwQKFuGt9QxOLd/4rboNp4n4FuEiS1FNxYuGbvLJlkTzjAF61ADcXcx8Q
7s/TKnFoeXL7AmqSKGwOXHTCwUwsAo40QrIEWLKMt3MH/Wsal7DsA+/q3DwJ5nOE
lJBrmzQfp1kWu239v/A6Aj09ViEdchwgSXG94Gz/fnzwnTn9TspXuhL01tDq/fnS
h6b9FhyOoRqf+B7BlchiU+unnL3gnF5nJP4jO2fFGUodXrroKGrNa/vYZuONVxlQ
v06rfO/9cx7o69/KVg0x4gFdUFuzn1BIDaAx+HtmYP14gmW9sGLKNOKlaFfCP0Bu
8y1g3vUvsPj+mJOGYRcL9mSomQF8uAwu+jvxdNDo+DcYUaYLZVXNHhskZ/PGrvKJ
p/HeOpyL7XK/9UkXW1SVWslFq77DjplZ9cm9whsDDQNY3c6dDRZONPQicC+pxl1P
iqfBZf/D4dbfJYPbPJYWTBeLFFItSsx1Y9nHXSuDQ+jhInUA0AOsZ5oBar1uT5Ps
efvVYFqCQ6NUj8e8bcTASsxcf9ac/hUIVtFZn4MHI6GTOIWX2rWkVsAz4dgEHLu4
UwimOBkse6hgTKEOdoWeEU/oPyJJp9T23/tjw0dQjrMRyAUpEF3x7IIsmOFpHVSd
7F6zdboUG3BsdYbSqCeuu8gUyKrtqT4aWiioXKqYO1pMp+Kuw9cXfSp0Uv4VjU3A
GxST3vj2npyWQYxsy1lE+D379FyqlVDLN6EpqbJuwOx76TFnvmERbKys1OuC/cio
KfcmRAeMmcQP5rzr85CBuZBYS7ziFnGnx9DpzNKfsMfPM0Wq7ybAICOI0TEGbqa/
6Je4yBZHE4Y/slJ7f/o5bK/ISR/XYEvhGhiIsVk27V1hPDNJOJViag494WwQa2bk
gTTWU+QaE3NSFMj/e3oT2l50qgZ7CcQHmS+xfYUePiQkhk4l5T/2uAQvsdkGeoMM
dY5lwtmXnUnrgS8C41H2EQO9SY4yGgmqNLcq0CyEt3SzpogWihXcJIKVzJ0/33ZF
Jlf84q+NFi5g5rfg5MmjWgfl+uqdJF70ddP14oJBJX4JkyvxEhkK/iwhr6CzjZI8
XlsDizec18eA14+I5Dop9u069JMAJqtApQafeDWf4rgbQDT/QpGnBA4iyFZdzxrO
pYhdRPu1+ULUcbs0dAaAiRy/63vDyVOoY54Q79J6juE0cVksw+dWo1lFewSizpWH
LZW8RwCmW5TSYRUMDlDs523M1+4ob5KXWJ19UtBEJeybhfyny62GwpOSQQ9Nb/Gj
7MJfZf4PHDIM+YNxrHTa3hjjziDTUg8hLQccR2/K4YFKoIyGL0Pi7rqonUsir5uv
AsDN6omqTwgeqUBEnBzI4CmG760xdJyQ7Ls7aAT4bZsAxNboW1TGGkWQoJekFYOi
t626NdKEUAe5z/YSxHZs3SKkv9Z/0k+FYprnpgQcORv9qk7lYmXoYQYPB+zWcHo6
MSJGVGr28AjHKW41AUIHggx354N625rwG475mCX41EWbayDRlcNnTKxnc0CNFoYL
Ls8T7yxo9C4fY7k8TiLFLFwpIxp0/aWe5I7bBH5QNemlb0fKQ9cDg+wltJO2O9AY
23l/m6IUGWl5VT1nAOHhKOnfcSyRx5+Z65hZeVmqdHVBCVzT13qwc9W+QwJ21FQp
na+rrTpuTgEm0QVs6uxXsVEmBU+LKxaSinPXAW0Zqd19Vw2sexGGnTgyT7GeGHAl
EVIQn0gzq87G5vkIpGJABW2GPTCwbLkHC+o3J4JIsM/XqM+ShHfDI92/fiYZ0JGU
xR/yiAWVslAtlB8SybC2qlOesd9aLS7HL8Eur3lMaH8sDZykdHVetE+edK9VHlSI
5NYznr7d+ax+6LsZHvP87hoFl/6hIlUiuOD8J8vH0UVz0KuhoWL9akJBvv/jcOw8
9SRT2MaGXVPcbpMCHyrNnGGE0fqot6i9c3VohexNrsQpNpD8E1d2MjlDQW1N49Hw
t6GzoA36zfqcxFUbZEsdtBw+neBaqSmO1UNO6znBw/hUsFjzRSQxkA/kW1uoAc4A
0IbSOR1uoHrzBdd5eap1Y4VEJMH5gcnVT9YubU1uQbmZVJUYPDLzoJIVOt48WzsW
Elqjw7hr/tobOHeh2cX6iVxxawOe0GB4P7nWkiDW7KL9SIiVwpXXo6j0ILTLyDJh
U+En5NL/C0I5GhEGWScCJLgehP/UXpN/2sbOBlVtmKzacjchJQavMjolvl4e4Tw0
ey+Os4xSVmBO/F9qZrlUbqwhATV5F9BvfyDjAiSKXLBdic92u8EoYulbYiRH1n/a
eNHY+31Lsfn13DEbf16XBsH+lLsXVXdIIVkDv2Pi7uC5lG4krJEVujEiYkCXwLIu
ticHhYMHja8WSZSlAdZOeMEjXhy2ojDJ2gUFq1M0kdC6OB/Negqiczr27ViV/ySE
hASehNm30JzryI7LuC1xh5dKzVTESamnsRoyzNaSJMnBJqeOglLwgVviA3mJYXyM
nntrhpt6gySd4wuJhvkJaBG/RDbkH2etfLerupDQXF6fd0kpawG6H4VCc5pi6PgR
6oP+6SSZKE3e5wEXR7WFlnzzh+iHE+suuP86DZkF6aLaNXzIMWdbkwloxR7x8i0A
Meoge/nI/fb6BQdEIu98DcpXct1KcGqSaCcTqzckNFpQ5c4QC9utlg48PuwKB9kC
no543dMCx+AMSELpjCd9nqAE3X374Zt8SMOaD11Qj/+F4HSaq11i40VFY9Hpimam
UKJmfZ1Se3XGpk7GxQdsBjxYnjj/kTaarum3j3Bl1s1HqH7iAm8pLRIANHXCjqM+
Bca7SPoxY/ERnu0A3thyIr/DuiMdwjSaRRMCZHPYD44EM2f1b0K+V3IIyEWVwn1p
b42kya6FyHl+5/iXpho7bS2XG4fhTdOr/FRqG/prydN6ZHrwj8nAp4tgXVLQfoEu
mmoT31AoJeoQmBvSIs4/T95p8Ms6G4XtI1YN4v8xbRA2nO7stGkrlt0nSVqxksnN
/qORwaDJqR07iKA5v4/TsoENa+h9Er192sre3aYhH2El8ghpVqXFken2FTY90qNg
3QbsjDRZAPOylZlwpzPHPNWBXUQI7bENi5IEUye13T25FJIVteZirlEvhEmIdq0Q
Nekmh2SAjuEJMt667TnyPVLPZUDhjTZRhGZ5vGUq8EVGNx4/m+wuLqFfwmuC9nDp
ZTlwtqtEfUDK7Y7HBKnuDhwUuRZa2kYMDbKauN4RpVFRH7g7MBYws0yK8Uw4f9jQ
7VWnotRw7EsXbjpdYGqsv1OueATgk2JeVGdUWNLw3imqWpLm1n9tgoF5yiLJKX2v
8VCUDdd6/cMvrg5ANQLt0JhGmowRNNTcaEGffALEOWwA2sH/RytDy4RTvP8piTnt
Newl3iCEZluPNLAbv3F08S1Eglt7ras5CVwSUa1ASvNh0CIAG+cvKLS0f7HpPBZN
hGWfNQBo54mvAq+trO0mG8D9QB01JvBqsdIydzbGP6qtMLuUC2sqW+k+5QxHu63E
b6ZnhV4pYIkEWWYJ6uzhnbJbXf1AoViSTD6ikA+XM1MBB7eQH2NaYJ9r6NxydHh/
pFw0UU1OcFFLtkXAqYhlMGK5nSftoRg/HUCjojM35OnmjyBLQJB0/Y87Wngjox1N
+ZGbSoJPUX+tsdYV1CgkEvskWf0JuijiBhE9C0VUCJRhCAxlyiO1cGURW3E+MG+0
UACYKuIB8MQMmbWaqNP1ClbfIN14cAtjxyPDdvLNsdb6d7/4zXPSgdJ3/YEXA5/b
D6KL+dPiShwkBGqTjzd+Eqm76v44/UNxfAuN0cs4AH1084pcAjAd01+HqCrPmUDy
fN1hwRNjtTbtNjF4M5jFtBr8pP2QxHzG8Vvdj1x57VWMUdUMImCx4+STkzC375ac
T/SrRQPX4vB2qBiCTziHiU85R+dtY4Gdg97YFW0ESOZlCYc7rCfbuc/v37kZRQ3j
3UR5O/rOcCYXMC/plXG5Mv4IuWyygGUTnUMHVJ/WABR6ZO4jWg8E9W1pRGTZxJcL
TIam4vCyVyaNw6qkDm4W9jpMa8UjRp4KdNozu/cQ4oT/ZxxnX05b6+krTtNaMXMP
a5ErK/YBG50o8dePk61U5UGN2H7VHnCwhiRXrP+i0J7nZmITIvZwSTHQ9+NXlGLk
iHgAxYI9/gM8WETFS1jsyB+5psUpAqnQMZPncByahdBKrNjoPrZbPHjvKQmyoql/
eQC5mEz9YyBlqeqUr+2o8yRB/3/6eZexqfOdt5GGFDMgzgwjsIkGojtDDFktTFnA
aZbzw7M6kCbl76ESqQqqWtRS61i2Hwe1J4rs60oFNpes6S0JtgPBQXFVlzbRH77w
/mCRVjU/DzRENygYwxU/Ww/cAcMLEo1GxlOMTg8nv8yEWf6ILxendOgfzLJJsnfc
U6eV8Q+N/7qeWr2sax4uWI8jvoUiZ5YvSSPtClSQ6qjeV8v9Sk2A1FDmxu+kDnLx
bNTTuDFSOsmKRpDU+a7tXFSigvG+onKkfO/s0rwVR7xCoHAyw8NBMeC4Jw59Rvl6
A4+7H4Q0DG9lbB+CxvK3/wVAIbA7iEOKJowu4W7EtDtdTWJQZwCHdbQZhnei7l8X
Gd2IU8cr+9jx6VFKRSp1BwTL/Echbf/VTsF94HwXZqxPGGZ186rJwynuSnmfKFIG
vA09pMiGQ4HWYNzRxGJ8WreGmcuVxJ7LrkKfCG/x8KJU2wE8ILojEsFc/PgxuLEk
q/+Fu/gzRsKy4RyNJmVZQ9YBx9CmAB7T7Rb4bNBQPsiHosDfOHG16y0ncjoXQp6F
wO/IyoOWbtSCx7mjcX6moOuH18aA56zILxQneoI027Ve+mJsotvHjI/+9Y0uDT5J
qCnMtA6Nd+6dGnDgPVQvs7/56SNfoaq5Haz0Jo2pIKX/A0As64czx2HBOrJW+9Fu
JxbgcywzTASVAu7YHNQTbhmBuBGwzUqd3fdUg7iuhJfrSMroSwhRww4sgidMK6Dq
i1S0xwVW8rgZ0EQklYIEUvp3T0Y4lcoi/NGe2RXZtCqsiHypxu7uzUc59b1Us8wi
dIVp7kPBT67dI2mwFdoyrAc67dMgeZiqui3LVrm/VtLAa9yKQOsdB6KCdig/Cur/
u1uH4koHpoplSU7oLcpGAQ6GH7S2I9AKcvab0u4pJEmLI3C9GcVflcH7i2+0U206
L/toaEacKkkvKUhCAvpF2VurwPIXR0VJmZ6iJuLj2LFZ90WHKF4Ubs2oA1Ymvxmj
w7R40y6OmdQqLVeU/yWMr6IDQIDo3Iopw5GozDcZGVDLS2BHMPoWnLVs4kurrBcH
9McWtCg9677hXTdhp4EPomne9uIEkxWq4dbpsBxxIEhdFL2lmVUhrtkWNzfpTtCg
X/KKOb6iRG9DhMbpLCvE9U01VU4caoKbE44S4PSAC0BNVSTuoHPkXCIH8S+P2b3S
RlPmHdfN9of/EOj3ieQwTHvVFFXRkkuwr3DQTzDNOUp+RIc7ayJuvjq/zCtWELNo
647mcrgngAWVkWzHnVPjoyC171R1v4onsFG8GeMRtSun+wVog7/EmpnTJymWHfbB
Cq7gvW8ATaoPwKIl+EFktVppo9kYbptD9tt57xWPFqHgG30Ns5ARQ6w2BBuMLmkd
rlk3bHoyN8JBl2xvArEF3ovn5ZwpOyqC7NOdfNMKoccy/6jiDuILnfu5tsc0/fEZ
j1uHwZlOTntb36OLwcdHvxKHzM2GbbCSi86AqiJZxPbGY37+XXyIo3p5Wuvkvfbg
/M71NjQt79teVVqz74CbyE2bQerybrRwwStJ+q9sJl9Gm1AaQcgWL2ZXbKH3Z/Rq
wNxEr0KNSPd88nr7y7rBiOkUp+hPUqfspHB7ozaOI2TeSFCRaMRBBgwO50zFlw7C
DBw1ddrBUneu2foXUnP1K1v7ZoX2J2ojeIiL2+7PIrfsujbyuCOilhDx3Vr8jP2T
ZUUdv5PnX1JsSZVecMo7rfDK+M1N+0btyKiBciy4c8yHQEoGKbIecMVpWGHJpDeN
CBEzrdOinTclkd+Gl5nWVD8mrOR9/tYS0fyDsEwQa7PGItaEAc0zGHGXf2ipwVt5
DNVLk8GfJFkmbrbRrROlos/BygLfm80bl5viAloiskEjqcB8O3F1cyTnMRqEpjqJ
3ApUs7543gKR/ZF8W2syB/QzCBG/buxCFV6MCsAmBTB/kZzxlDR1cbNn+WGHtxto
UQausZyUi7QCVI29GXq/Wn2o8i9hGSVt8d40PffIMSUYCKAV+FoQZwvEM16B5ZQD
5MDZ4sDkKiP8EkzBZeFOoPEb0tJDDPcp1IWjfYY7R6aoKkMdBe2zSbb5me6pEyTe
jS2cBFq3rss83SQdaAAWVU00LjKLC4fE+aQtaJj9GwzssoWzj58ciTtPfSK08LgV
7WIS9BM5Z9FX2Y+77e6kwO3xFfGzismVEzdcGu5mB0FWrCFzuCwsrsS+jtlxD9y3
mHMnTkWu6D/q2tX1f+LYbrFCB37hetwgjuWqnE/iTuOY0EQv5IUbJN86eprTdlFe
D5P218ivuZCEc4oBb6jpW4bAKAvDNgRhv8RNSZB2Ta4gTa+UzANnJVn4ElPXv38d
mXG+RLKCb9XfUjT5cahCLcj8iTDYanD0DIqU39bAZdpbUT/mLMnXeK6LfVib/ngW
aO5u+IMDsP6Bf8v373uxU7612AmGhlK435u6RkIwFb1zy0GGruQ4nFglkEO6fVgQ
H+3nl93DGMiJjaLVXG0c1PYNsbAWgT73ecTrwK3gDtRy/gounK6iBEpHqxlpRoic
TQidjrBlWLrjMrOXIlS1RA62+Mv6gdM/ERP2oxnK7HW5ovmq6Q0VuPjto4lwNnL2
rYuLtYuMFt5SLXRV32yVFYUt4ImtcGQpRnS1P/hq+So9O3v9XdIv338e87MzFT9H
QKzuYHhaoP+Z405ugb9xsPHWkhQLu3BOqUief7+BKAAUTEOxjSGAXKgg8rHtQIfb
LY6mcPmwW3is4S63jgxr/HeVhMlzh1eSdm4pyNQm6Yj4uEsLe8cxMiA71t3VGhRX
wmd9CeFR3uLYAluWkqlmUwxwMq7IoZZi6INPPnO7cC3saVRJmBIPlFJQEbeq4EL3
yRdIdv02ky5nr/3UrGnCwnMJcmG5ofs572KAxwGn3RMhlShCLTgybH62jKUV58Ob
45+q83Obvjfx6kNO8/HtYeFexmI4yUBRNGQ5wkt1KLUlv3bxqL2IkEOOPOdGXUjx
HnzU6X7OKjW97G/NTHFUJR0QB+bjRa5CaISTf6IGqCnMYReqDva1fBryvpSDc/F3
3LfMksrlb9nb0GEfnmRcROI2pI1rCw/29seL4CabKPjRPYJFjOQ1XNTVYYYnBeE1
mO4ceKFHr/wXG9kW8m+Bo3CQDqvrcsICnZjPigoWPF38WvAalMT/daVj2TicrEgF
8+XD6i3c4fveL0A7jJoNGySM2ydTdFRiXeqEk1HoSFkSiSOL55ni8Lwi+6qjpxp9
OYw7aVIMqhLtcZ1NCUVQczQ6hnU1D5wxyYO/0qhf87syxi97vNiuGjt8cjT8izHn
msp4UqUQdFC966PG5l7wqSi2/s+vS2p0Y4j20m7YAkq8QpigzRfGR9nDfm3eLeRH
fFEYiblYZnukSt4aqGmr3JcWOGDSJKv+nPW3LYq2GSBV48/xIWaLntN+sz5UiTJA
nIKH5v0i8T3BuPrXNlcdS1oRrT5ic2sU6C7Kcj+dyhu+nT4eFR4m8/U6jEsaDQqd
V3DzgsH4D1kyq5wb/75Uhhhiusb0KLEwyayioi0DqkqjDMKIVYC9+I8sSMswDEdb
mntiyMuqjbmrXLS0HR8DP2B9pAsBzsKQCePlSbKPzK+QPo8dvtsJdKnw0INcCYXc
LeYRj0w3cpupr2G2Uhmy8TyrnhiHlFGwbC8jVb2ezL61hIJGM0qZOy9dlR6HFCt9
pUzOq9F5/hME4FkqVxLqVg0ciwAUke4OG5LgwZHisfZliPojbJWKWhfoQRAtac3X
eyvRIB319htyP2wTflsjj8tK+OIdex5mUEXDKysq1BTaK4UHZJD6WDhP0Z1PaIqx
p6v/muQWlDdL4oth/8gaLm6s9rB+6yXxa6KivlMGd1Qyq3QhwuYqHGOPJI/Dxh5L
m8eME/KJPtdgjgl1ET98CRfsOaGaPEN2r8DmFvtfMymOYauhzj/dgM8tIMoo0IdL
sTcVj45vU65TqIJcUoS9/aA2FkUiQ6CM239olxvY1x+PNkbTdraHqn9EXzxamtVz
mbuCWEVSmwANt0gdheZRM1WbhgrTIbQp6ZXQmeVn8gqt2wuQhuydll8CpgIlKiKM
0FoYzbr+vG4wgNNIkQywjVGxUgT9nEtTi+LN/kK2n8KYD/Vp27vOsDhrgbIZu3Hl
/nfwC7tzVFQvfU43kUNELsAWrW44SrxSYMnqFjAsv/IJS0tOM8WPin423oa/dGrX
fE+HaVvYnZXve0mB+xwzi63MHf9LZFgZUpNBWLsvA19zY08lMeNp9cGjw6+0aIoV
lx18nLSgkxRhaPlY2FXC41yMvrgdIQpP5TNZWP/DjCTveJeY0CCMab3EJ/rkJkvh
WGJz1ptMH0wWrVy2GFdLKLaTT0XzU35I+3tk+yZJ58QYTkck00V7Qlk1feDPt9KO
yzmHSeXczC0uS5WlwGmPht+kHZWZdAr9EMo41AQnX7o4lYE0Qw7nx1K6Rf5725Av
IrtbAcZrAWAidQUFN06+VUv1Eb2Ig9kc3CJSwio1F/XmGrHgw3jyl0xtoXCsxNJh
BKH0YlLgNMSJPtMyJ5qFnaxMEXQhWrjkJ5glfOtlUs9D/WGA5gW4kZMst3FUX4+T
hbpuXVhBgtIfyo+MhpwYkfKrKyAE4CcquwSYoB0POTA+8lSiPBhPKCkwIF+tovjU
O7kob2aPnFpDaqQIr0vhHzKhJ/XoAbj8O55KvzzOUwx9qZlD/B0osjQYRAZ2EEw0
hd/g5Z78H3vBmAHBJIJRWcftW7Gz2do8hgx9DioU+gI8jEx1cpbsDorh9mxuVhxn
oAQCFCdx2H+lFtge4o9/q3fEtPx8yCqsv40Bohm8L2Kfcwx1l51OZMb8bbJeZVsp
LxIlEUuhaWCmrARte0WpnYGz1blwqR5ItsjdhUJh4lGrH4uiumWkg6T5bh7qeZhI
GnEY8f+RByjQW4Lg1c6s8Ehu1xDP8fgYPTZaVLbozbbGgpK8dIj6GgC/3KWrgCuK
AtPvDICERtXbJkUMjWADq74rtZC/KqgAqhTCmjxfS7o9E6kJpn20QrmyAk6h+IMr
JKjm9/tf4sAfv8LjmCa5Cm8Y1tIze37SxPmnPq3aWgTc4ShEsIGHX5djgF6esgH3
yCydzxA+cortfHdanck9Slym03glcHthaRCLNykdKaPRmZosfHZsFKEeOo13/gM+
h7IHUICtrppG3F1RpykpUJGN1AxPyVy6DGVTreW+pySrCy9NjaD2ZeZMqgx3iePZ
v8neTF6EtrgjK950Rdqx1qKtp4semtw/q4oZp6baPuI25dtwHvgjKMm6FKr9NKJp
5K5JSMLUHPNyxOrEr4uQO7xVyw18uw09zyVOb65wLNxLxpWomLfDEH1KPsQP25kU
R98LJOQNx69+VbOeD8jPXqa/hM3j5NbEVX96krdLe8wZz3kl1zqUzRRuv1ox91YE
yZ1NbrzYialdMpgp6a2tWw8T7Hzvoj6Y4Vh3FuK20cCM9ESDjlpjTieelQDOxnBW
McuI8/ve/SRAXoOG1OLTFo4BFBnEuafifpiytQBRiV64AIAygsxkDP37KIIY9vST
4pqI8iC+ouEJogqcqoru99HZhRCaDgnoDzCAbcEL55y2AELmy0UkVassjV01PBv3
9o93CvuHi6ZEmtP1kJeh4/otSuv36yzMElvlK3O9Dk+LXUVcJV/13rotYKe06h0K
3HU+/zBQ26oYMr/0zos9l6FJHprhmKFeN39GKwNOxqWfZc33hZ4Fdv8W2jkOWYe0
vv5KVZDlIM43haDbNpvkL3qpuC6IkPtxddR2zyJYx5wjBzIkc/fyOu9oWGgkLRrT
ndGEjpook3rH4+bmYxqbo8QkyEcGmaLz52P3z8DOkY10zOJPbvimwEv095+aeZ2l
Vd0eRujoKOaejyFhogoI0oayJdKpnGaio9J0czrma3iJPlCzhI/KankVTF4AvZT3
NjY8SzlubjWItBQYuNKfRTto+1JbGXSiKPbVJkC8+ghWO0EUADILjCJzcaBxa/hT
kejfTASOZRBxW+7fA+w6Bq74B+Gl3U6+jkbz/pqCXg+a3WbcYAFeI/syo0Q6weGt
OsNDEYQiC2Tp78e5izT4i2NsTdQp6tWH9CErbEdQKp79C9/wvsqOcIbOA7grkd0N
BORtM24S8Lipd2fy8a2EiLfN8UH4mjEg26B7JbGNk+7Z+AYDg7yfdMbci2QJ9GT3
mfZSfXppiIY9BJRRTb6uCc5SH7LpURKEjpJ0WDNkG1Z5lJz8X4q5Mxd9M3pf5v5z
eJ/CLRkhAANk5ScBSc1ddRS3oUxTKKuU18mr3AeTdNczJ2HVTE6owgDi4u130R4s
UoU1Hcs+TXn9OluopXSEPEAl1qSMSwD6Bca72yVtHh8RT6pkLZUeoNzMU5jbAlf6
7pi/25eGTwKX/JXbj/Y5+ToQWo7kuIKuGsUnXfQdOmfZ+8iBRyhSEDp3v1oxiQuK
faYpwOHJHPBYbWXBJbsSMBjcbx08jErSFzrV9RbWVFhmFf3UsD+BjAiwMa3LMX5C
kB5swvEKrJbceQgWRcwQg1/eh7zDsSJY+wNUo9jC2G5waPrdf8zPtDqZYMcv34WT
RCt9sNEibLoij3fkG3Kq95DTCR5MGhxTaa6Gb5i0FiP5XLTOCWYqy3UhOmNFdspI
+34WQid4zNUzHOqDbVk0jQ05Cm/yNpLd/lRUzqDh1iiWcZvE5jrpHp7J+5YV+lUi
4BxUc5HdLb+TIyPJ+ifC7sfgx/4h68TTAknhxfZ/C/jIcXhjbxKKK3w6FejOoVg5
hWoCFpVQuVtWN51VRkgTmpcRP8SPRZIb63CBK3S56C7EmK7XeJEBAffe22B7GL8B
bFfU8hJnI486qhVyJtqCx4TOKPvXvUkJW/6uHDgwRwJJSNkMBFIt3GnjBQKVaS/I
+m2nLz2E5xg5dR7yaodwCBd7XmIW/rMCkxYn2JXu9iXvfQ54iYxYQd/zymPP38LO
Bpn8fFlhWgopKR8IDuokZ5uUR4NZe/sHj3SZoiDJsSyJIXb+YxoyLgvz4e3i6ex/
NNPOXHwOm04Y0e1QyPGEXj6UOiOsfQp3Q4KJuiRk408leGf39zQu4ErostZOaV0Z
jK9ZCJUat1dgutnpUr69EhgxiLzcG2wgYLbNfXp+h3WS7LzhlB19+3bsVBPLvcEl
7Wz3PYR77SQpCBQ/+Y97v4NycEFZJ95qndsdGGX23T308z/CfttWWqkIoo24pJOd
Ahfngol4MVAnsEbT4Lzu0+uOTGjNTXB29YH0AW1QdkKTkYmMGQ18yWVjW5rVzMc5
F57jypKBcxZF9q0iyx6Ls0B+bG9UE+71YLa7wP8tOq0DQoiVjbvxopS121eoqRX4
ChM5VhwLs8CzRdO3Z/ZIDs94Z6xwWsfC1Sg8V1YowliFYCYitzv/vMMVjWLY6ob8
GOWUMDIdh2bS0C8kbG3Odd5JOXlDYBMxK57lyNB3fvoHifY4H94lFJGzes+zCtOJ
NyyjRfycrC0R5QPe+eAjJBMWBW4nvMq0kPyDNXHaWhd2W5BWGSQVYzSAZWQAkNhZ
XsdfpSE3Gje8/uA5KxjeZ/cdvY3O4TF3S1vr8HYMQ70v8tR8vIkM7UayS8Qqhi9g
+vkL71ylEnzJpo3tV6whoeuwBRyiQaKD1d+BMYRyuk7FVDLZaXp5QcK4YNw3OEDe
GhmEIcvf5csopCH3K1F82MJBZ+xfz4vRWrAN+y448+dUwMmlS/WVTRKrikucqbYr
h5Hc08qyBzxGDo7Ud++KAAb9wYetpziDTOTPZTbFXruXc+2MY8utLgOAfw0qDh99
ni0x1G1idIHEnhY3yz4rrYldB5E38Y8j+3FxddysKvT7lCjKo96tHXbhCHaa24xN
C+XIb7IYtVGvy56a/tKS9+cjqkd0lRl4tP3/BuJafvk9PMGNRrhAk/0j2qRRn8pa
IBKYrJQkJfG3oKamMlrJpdMvJ//h3aQzG9WpsOrrfWXxk5BE8JP/LWWP1G8w6Ler
cTnPda6JHxb1HH0Ab6uaqWQwiIsTzeNBP1zSzPFB12rBzWezuCLQRp+a433yh+4L
dq1eEbEZFINYClBG3toLkUzyeAynBDjGCmkD4ppq34pM7Xdy64GZt+4HrrKPZs67
lBo83NEnqob4Adv4aERZpGQYVSzVaLszRXLRfGSC/W9QFe40Dwd0W8W46wiDXNyd
n9mjEQNvEGiII7tUqMPEXz7wsaoYbes9uvI300xjulcGSu9SW2DxVK7eMYlhd/sy
SJNqHaU4uKEiOSOpoYJZmHws14Tu9xIOtQXxtexw1pZXXJ/ZAXWOyLWZx8wRl81O
ucVyCSCz0wKk8Yg9TY6NO77IpU3T1p34Pdb3Jr+zyoF5Q6BjeIkRKKaKSLaSkp/f
uNQZHhd9vBTz/Y0HOafHBpJv6Ta6txoAZY35j7UsmohlsCrCfDCZjc2TKRAvKCts
2XTAk6hP++zKPQb907mfFgGMmAYcp5kRPxkRgKAlyCATyqTUyDejPCK9iUwdO/AY
VrQ/kF7bilQd3okBSNixR9emtYtGqNS4ulHfwcxycwLY9I/U8slfsGGwd1LvvEc4
DGAt79VKoRv+QJNcCxIBLVH4OWL1WC3nGVJIx2cJJFlMkelh2v2rvM2fJ4fI47Gm
vL0FYeO6TsYiQzpJ8kAR62NahYmNoAyMtaZbTTOdnzQt+/2FHhmFv8uwjdHjHPgJ
ICyUPFyfPA5GBJq1/iaICam0Y8SMPe7lm5xa3zCPN9GWO61GmZd9fu1bgy3PxD6e
vd4xxzWCxdNLONZB2dbIwL2+cpN4EPoZrauEWyTIAQ4n40JvDJi5+qOmaT7gKuZs
B9W61oF9NE+5qg3y/LYRLFELyOEqkrZaSvy/zqx3Bcp1Du2TYrKSHp1/FMrhzuT0
VvFqfIc9DYolQUaI70j/Y46bNRbc5xrThyAsU1MzFGT2ziz2ZS3M2lUMJPYEx2ji
qNZDBMDMhjapr4x40Mazt3MivNczXqBAf4UrJLk2BpTxgf6RIvNPi/qJlsmWnQys
+yUvwbyT8o7J8bq/yzFKgD4k7s4kuFXQl6QH3vRD4JoGhOOem82qiqP7aJ8A2XxQ
2UtfID3k6rSvh8aUiBPddtHEH7EE7BGseJpMU7u/QcDgtkGFKhmbu1gX7dkflyvX
EkQ6jIcfz/KDerbcYXCymO1divH06lwY3uakdDEOWAeezB+icPtvp/mwfnP0OSgc
Z0kxr/zybirDL53rAw/LoKm8Hg7P6tkG5/08FhGtflEwzj6AJT8KdGMq0KXM+c+x
jQhSK/8C/d2lJ5eMYLVAJbhjA4k+iKVnqbW6EjsWUsEG4O5gP0hhP4lfccFBfANK
AQqjh1VUzuMet031QVdVjw5/VtT/boeYDhHWBGw5plYDvMqoTp12sp3hrG1o7u8U
5f8svD0DS/vr8I+in3HxyN4trgSRBDokmw2PHmWdZe4ZbJevgAUBHNmtUJd7IcEr
eMKKtLMB688kzmGQD7f5P3ovtcLuCsuY3jLw/KMikmFiF80IRYprCa9MlGwud0Ky
G84BKlPPr/iS9UlKyLWAIwdvyqk753bLTCywTiRX6BR0qNjfxHPJI0+68an71ajx
tq+/8LZtsWxExOekar90hEdsfDhaPwVGT8WDiN0Dk74U3Plwiy/S6pnPVX+uMqsk
AhXe6xwgpyeul2opQljREOniK+3PK9D4t9gqhe4QMK80ZFSHVhtCrozdQuqrglmx
QsyAk1jK1c5Vn7HdByK82O/uW/BLCVO/o+6nv/FogG9BjUf+nIvRW9rS+T64Yfxs
CveuVRHbOvO3kAVkjPEDSVG0UAT0rlh68w2teBSkIlORk/tvpwtiSNntqOdJ7E23
1j0wlI1OhmIepu406cvoIG44gFoh4hc+0Y7Xk3igJKfjYTQ2F/tgsDlD1yJEM+Pn
foDw94MrORuIUeJsh0mNNYJLYfn9HAQbh66L0Xi0Pd19UCaSfkz6pZQJShNuITBA
NxhTOzzSg1/4Fee7cAnQWepnB6N+76IhEM7Z0bv+mv27fBnha3XzQpaunpk6iFH3
2TCJG7aTM86K2cYiLMiI+ot9MX7lr9xPlq2aqALo0LCoLC2itRK0PtNmGERsXsUt
XcxHbDVeRLLKidc7vOTtcpE5ktaWFpnKUF7jEKgw6JjXYsslkatgqooRxm/JA4BS
laL/EuWVTStG9WQyCKMKEdGip1gs7VlRvKH9RS+gCWE1OgEstYQ+5uA0mzOzQ4LO
OZkE5jM2qqGX4XEJYiZwgE8842kPufq59vGAQaGud4TawKj0pBNncgU85iGATPAV
WjBgGq3rf5MaKP1wPfbnZ1PH9MgZyJoSLy3ZH04iix1EfDRdXuHYTOwsZCa4S4WV
c4YmbI2KKgFu/e0XNhht+upBeDySx/MiJDQsDbHYQ0eLMyJL7aQDB00sE285YZNU
KxIlKZr549NO61tKzVxxo6mynTek0YJ0rPl8W36ehIehedlAWeYBf+CaGi7UIxa5
b0VXReVV0ruH9a9CmjSPTnjfzSRRsxd5M14Mo8oN+QKMIJ+btElqROc3RmmIsNb4
ao0Q2kegjNLz5CU00pHHB966KufqLQDsuG9JwTx9hpDwiOooQMmPQfLi3GkHTPNv
uerdxZHR/C/KgEypSRp1rrSvGFHu7FVs6+8sZPfzA5zRw4cA5KWCmwL3eoKb0zZf
kWNDHFhAd4d2AIy/+vAL1cLUBkYD51lAMYiEYEpYOahwk8JwVnLIQtIa06l2syDd
qDkBJ5nZfwqIaiaEKWB/uxP2CU8Hbs16R68kWq75L3keS6vIj9M8J/te5mg1XCk5
SYPgS7sR9GqkDG97zZo+1KbR8DLft3jpXBmH5zD+YyKAos4oEN15f1Fw39TZMkEf
9I9NJjiHyKq2y2GqzqAtCgTUPgQ3m+hSX7jZJCAvrslShpHnQVyF8gC7upTOZfyl
1VVVFZ0CI7+uUDTs9UogUYhx+Bk7sE7t9dOidfCPru9SSctcZBUnDyAwBz3BJMVD
s7tVDLH/C/qJsDMtQ0esSjDM0g1LlQ3t1KAn7Yuc+8h+RHXKw1TJpGPQmL2FoJib
CiasMn47bMx1EnWcZNTPiSbxS6PNwanf0YZmvAeGu0FawWoXTevX96ieDT8ZYChh
liwcuK2AN3++5JuZjPEEOLGFtEFI2A2StqE2ExqKTsXPvmbEXZLPKvntsnu5HYjP
TVcB9usEifpOZNHJZZJ+P5LL4tYt4mHRuc7RawIdeJx8mhAlPcySPvYY5YDacfoC
amfU+YXbogTuan8lAcNOve0D6ZDCVKYkmD+AXqNEzsx98jYGIepsEIjVGqo7gZTJ
0zAqwpErYSNq2U1HoVe6Z16bF8qcOIG1qnabXENmY530/X5zWx4QT23kdWqkDuoZ
s8lL+Z93mdFZLk7sCzTe73fxr27HPyhI4yAXORyStKLGQmlioj/JTtXy3Cld+RdT
bCDeiCQGO5kIrsWwtGADP4btgjUQyIpDjeHu+XuyEQoj88jmtpMzMii0Epng2Z6r
0JUBkaFUlknPW1y/m8gnnAiQ3I8VeJpFre09Wnz55rMnOk5bmEqhCJu8T75iyUNp
P9XUXItue9fDSrjGsi1yoR7p1HA2wWBDPohQyJzFowPgTGvzfjW5VCiDyaJEMfTm
bqCdYgY6tErKug9pjlwUkAShWqgbSQwOhz0KO00JR98lXvGKqVSivCiIKuV87Cjz
iwkWXLb1ywbY4GRZhXOk8fD5sffWZE2J5gnT3IfYkCrL73gbrhz68Yol0nezx5J5
+bRJfbXeXtw6bdvnMizdUsYlWVA95Kegxog4RhiTo8KwxMmUuvhkLzaFbHr/c/JU
11aDRMj4bue4GjBgqRbjXxNjeIDncoXBJjbVKqAI+V+DYx1HAlifuknlnDC1ymtR
TfkhyK5E9O0HAPDyLqzEOLA9bTVmTRGFmUMd34NUfEzJeJRacq/OWCT8hXlcHU9+
Av9I6EKI+KuDL93K4zeP0TJ/V043FwoOwFiNjJM3PEybGzmSB7TOVeDVdfXZGGwX
GWeCgZIIAYfr0IfHWbODOU0LH3V2GBA6GZTE96AWagPciUfzBPa8m8/kH3rfVlF/
bekBWn0wbubayDWk/rEDA0MOqjXCLnzXytJcDc/Vi9C/OmsJVUPurAAdeTDYJEs4
AnGmuY2CY4W+mhcc1xPNCkt81Y5sG6rugc4cNiM+ne8tMBwDeNnBRwPxYOvIy+x2
Ji74d08SCLYIRdpevbXxx7cjkhcPd8cnoeCftaUQ2HJ1pvTVngUqw89qdxY+2lj7
I/6IEThaPAddV9VEvq//l4fdMGAglhYAb9kjNszfC3vvGD93oHkCXE+nQGpovoFt
C9ggcgiVkMS+gOiz6hB5nF1Bt7JtsO8HaaDy9fx/DxKVDYEo6o9pVPMbtRQ2P7Ei
dKjfOzGJmG0YBVP2P1Z6Jfxj7uVBi5T2N14Dlz35eUlVif8GcHf8mMB4+Qgn0OID
Z3bqceihu74UJmUA4pb0Cv1ch6sxwNs512PKdXySaW/cWH3FGfNGS0Hp4JTWn2R/
DCTmkRnJeSbmHX0CVsThC/oS/NymRn3tUOdbyplRBhqBBm20gjnn5a1TxGJ6OgcE
TLSq92ZTZxMlD0kAdu52/n+Z6NaLfcGUxesKSBsg0i5M3evi0sqOYbpaBNBgGwOD
AhVjbT5/Aup/dkSeueYM3L03e6Z4xZntKFznuBlnnVW596/F7oPC2X5eQNy18oKa
Gz9CzXVApfpnTZfpWzupigPBeugDwD5UuXfor+UASr/WsqJmgqyDjgnZRtv20H4+
tbpIg7NsX/De/E1GqaPUo8mzNCNVElCfO96ysRPiXDOvbBuY4Y6pjQniLk5YgpKf
A08Ey8NUlbo5z1OpRiu9KOWMQwvDr/aBf8ZcICuzwwzz/FXErRo4y/APBkuPAfzX
NsYxd3SzudEgX6sFKgi1qY3W+OugPRKUoIThDU9X50OgRdY0XbM+ACFqIthKxiTr
wYUp+YvyFcCHes2yQJ3Slj580CLuMtW5t9CUD8uw3mKGVEgpTCA6ZvW/A4/Yu3In
BxT4e+yN2lvznGR2s+HeZBgQDRotl0cB7jPxuHe3eru8T9nZ2GX46ra7mPwbbBeB
Pj+Xh2m3WIyDtrtkfNyjyOA2NHN3Go6bzlXEbYXE7RoKCd6R2hlRQKcQxVFgZoNj
93tVDbATjFje1tr6HewWVfJKq0Zp0VWGaYBJl2m+JkQtUilFPF1aQqJpUih9PQ7P
Qoq6ZOdG4uYew5SDjw3sFy/YWIhpDvhyamikgAthKpkquBIE+OBh2DiqvcmxEMsG
Qy+D1KyRFpOqiiIkGrHY7qSfaprzkCE2ioB5FdkPgLfuDscRPk67nADwmMXQeguw
ThmTS1Eb4pVEvvAQWza2H68byxUDDKdo2+zJhnT0zp0nLWDIkve1YSSGv6F1Oftm
20Uq62u965KKEtbYAr56wWYFMlohETDnqU7YcqaQtgPqPU5b1OLK1k0qQGMa/GL4
4FYqC2QzIO0Mb6lM5gSm3f+OzOc7htcO/Q5wS3LNCXgrgHJjJSwlNv+MmKN+3tn5
x2560kYW8NyOSMYc8wzMDE5ocqOO9QZ18rNY0KsWgVSzuRu3LppQk+cy9PPqzTsS
dv1bUSeyQRnPA48DsOIV/OPphmveJmanB/r7buax8x4w1qf8YXEI9cGM/E+rhMo/
NIGEvqyEIN7G5YTQRzb6pXZG0UIIQL/ePNqh9DdZPisPw2LzstrsA2epIY6wEDHF
Z7BHWP3tNEf/0736qCHvm4oERAlQ4ztdhXwzZveyNIF4J8bbRjDsMThao2xqWe8A
wbdUBjsXyeDxYmOXdYqTqqTEXyRV8DWX1ZKOZ1QIiEj/M46jTQhzuiUY/madNMw2
d7aBaGkJ/x3viPEpMkN2H4Oe8MVjWETOe8u2VhJjySp61CezkQ0IspOF85CkYFuM
jmzlLbHFJGksc0Vr0QYq89gDQrbt3KOClc5BuvQdcrqLBSPGSMomvLU71zYfxy25
LpzGo4Ilv3ULcjhiC4loeTZYd/sv10CHrurKIbnmtozT5xJoYjJooQj1ALcV0RiD
MoSFcyhUwNrnRsiU+N4byhciIjCoDtD1CNmjq7rvdQV0k1wXNw5bTQbcjol6sM8K
cYjx58OP0qFsIoQUqYNV/gJzcOsf5dWaBrNxPvg/JS72CvPPx8YtSPgqnolV8NgE
RP8WmfpsD59JucR8DbfCYN7wughQ/IcQeATz4Jp7Sc88qHNBIaftnwCMf2/w0yGH
XPMFbauMSSgqRBeh2A4uZQw2+TR/hp+3/71fsW05A+UszxyIlSIRaUt2hzT7hH6n
+ctRjvirJ+C17Jpef+RwPcRIzQ0CkfBLGrwczHd0Kf+IUJ2zjNg8P9Qr7AJldd6x
7wNw8ytwH5U1dxRfNUvNy5w+gUQS8UiMX3f2Mxrbpxk3c3gUUE6bUSMm7+7dtcbd
rjdaA0fzaUY9T9Z+5o7wvxISz1k/QljosQwNYnKu9tggTOBVK0PkV3trHf+IUiJy
qIfdqOiLjI2mkYWwI+kgGUi4r0E/B7eFp1QcHYsxIuA7bR/gHtfYwPRn3UZqisOz
NZ9rSSJXNVT4pp8pHFCUJRT935tOkmMF2li1v1pwRSoRy+4SUYZAq8/hnoX8LpPH
v2bqxYNWwr3ITOvyUjzebhowUkgxDYAhRjegbFvWow83+cfpsQWWMfojH2lTMzMM
RbeNZNrfB3/UdcfAqgQWgcmIp7v6TwW2ppNbyajQk0mkqDiTnzYxila3ZepFGY+F
X2xwuyex/KZ7aYrNkFOBGKv05KeYRnsACWqAPz6yAkygO9b9GPXEXhuIeWMj9ciZ
hAz5yLLei47yWq0wsb8t5zLAvZ/jk6LUhlM2Cy/OLeVjUG/CfI4QmI8cKydCHND6
ceVFlQDJJmorbaQghjpA+0mc22TmEYALANAYsy7rYjCOreWBJDF8fWdYKNHa0dhT
1HbozN07TiedEppP2uzF9zGOIWpzEZyBmXVfc8/Ps47PEXKG8VASk9DWhLf2mMTK
QFi8JMxqLGU0PmWa1daEcSAjzaPUpmxfGQ1k2wm5ybWVWpU+CPwp2fann3j3CEN7
2H3TB6rhiAYSQJaDulkNRjDOKg1QnMv9sGezvOB3RtyzZ87lx5D0KVB2cBEZ1b2V
l8gh/6HRUosaC2uDVOZLNa7MwMPSubVae+FBvqXCI1/uAP2ne8y2xWlDwswmjOIb
OwPNfxOEbOFRCMBv5RzyVEq+mkGvYXTzlM9VWPkDHyJXhpFgZcsRzSDBU2sHdf3R
B/KT5uawAWahabr+QuCls9Jamdj/wQAEDXWnYXXBoCAcs7103QwGQ1glq7EWLAVs
NJfggffea+4jlC3t0L/oqQwiimmCm8AH2UOASjuMD7vl7Z+FEf9CQPSYYvu4LuQR
fBpRMuuuL0z49jA6hIIZLH3PMQ7RrNDnV4WMjxBW73786vOZeL73K+IxOLq9Zo6k
2mvHe45yW3b+GnotaJ0WyH4AnlxvyAMwyCz0oREeJK+RV3yVZXey81NO4OUhbScP
6uh+bkUKteOincabUoYI1CuCOv47f8FzXTvmr0W+UcF77hbiJXe6eAmRhnRPZ4Bh
kDsQvdTVzeMHOWTpsdVVvOM8cq6b8LKM39VyXi23n3RNBbyMyQ80SbV9bXi+xZEj
Bya4rbPWmu/PcTlIW2VbB4bjFIONa3rNZBb3TOwTiDLRhPpu7tVFVdM3mZr1Vl6Q
nYC+D4U6UpBd+SMoE6jppx6YaxbulAnQnTkK4qRLQZnN0Qm81r1KL64gTImG2qwS
ShEf9ylZSMdLc+Y2tAJrN+calR6ZvPg0uc64omS32P4f6PI8GptjxwHQ4HGRqzCr
hu8VnIACPn3yM90j/ppqnoyLii0VzR2di3EgZFfNsSefog5QOXOTP3HzbA3ucbzR
wbltRpxs8hgWRpLJwR9qYnLTyvkRaADqbkSkReb5p58p6EaUhvvsguS5uwA6Rmxa
Pd00TDrTztBxfTI2UgAONq6tGQYTP+L2dQsKfXLsUSmbmyaY6IdELCSJbNDERaU+
Eo+bRxYCorca7FyUrKOXdXUKQ5VE/GkAHFFD/GEL5KCKkVUeNPO3KnqLNth5jGSb
LDzINf5S70vN2vdgb5ZAH9WQVdJe1LXfHQNsrxhwsJRXeCNfGDiPdAvLGEUm6u4B
HhG8QV6jE+/nmvkzp/Hh17Yu5UmvRT8HhNdxHk3uyiIQDOibg1V5JdfOWkn5l2G8
b1v9x8Yyj3XXUBv2dxGsKIfuXCUl5gLkFlzbUX6NMDMI0Oor1rKMEkiTux6984ui
XRLGszSWKcbaTh8LNLSBh0c16rkd7KbXF7NiICZot/4r+YNC7UZr5dxQTEDWylft
XYlnmhMEtPcD++iS23i6PF3i116wt8VrJFFHBIprzE9Jdo5Hr5Aox2q7U1es9KRD
lT1QQ+lM0BtXzWeRQZ23bVUnQzOXAqz6bPfWQVysaRVsYWmFMQ+x59IXEwd9mwL6
+SfRMh+wGmGn113KqR2zk0/vgnSxoTvnf38c+t+ZAP+k878GsmS8o/1NWBW+JrEh
S2x3gO5r2xYdLGT22CeMJZVq8WZJEfbythFu67QrMpsJuV9y95xz/p6jxr0YSoZC
/BHtQIwG5ZfKpdGnEKNo4GWOTix6DRgeUNWXD3nKixN3sFlBpEONgPHD0l1fVGWT
IUstM+j7Hk0pXjbLTGb8bXb2yCIDpBPA17WP7zgx4ZwZmlYKxAOIQOzNr0R+dbxU
mFlgXHuyjI7lqCy5cvYHH3KVlyTFlRACfUYzznwbr2y94hInSWL+pExLV2LfoRL0
DzFUbrV+y/QrX+Ojez4kz47QP7B7+4GEcfLP0JxZpkfSdmsviqEILFznYodjLN2G
WZ0vOj2b2YvqgBDfSOJvP6je8uPGtA2igHC4Q6FpyWI6eWpy6SHPuu+M6b57oqwI
X8xiP/B7CAZs1pCXhFEUb3n040dtFx7Q7w6rKAsHL9EWdI6ZdCuIVQQKMS0CCjRI
LLjKf7IMVejJkUXMGqwmk8iqfJ3DY8RQOSNJkQnmlnoyr7SM2jeTqqsOKR7op8nA
ZEFLmwTK3kZ1NUZXvxJZCvCiK4xgDwvi/dI9XpA8wOYp378obsxFQB37ItwtGYBu
i+iHtKmC3aWKKCZT5EH7SdTZS36gwArwq0gBNb6eJ/tyk8fZ3TegNOo2GaIHDrbu
ytzEu3PbwHa7U/0XfY216DPJW8WIYiW46QSQqV3hdRLm4lroaCc/Gi3hpnNmtwnU
aHuDZeIGALfE0EyeCV+ugc6s20F0xLalyoXkDFml4AXHVs3/SmXArTOyZ9LRbTDi
zGrR9DhJYNqE60YYBVzzwI+r5fuO67cqtSlAsIfF7T1aPVpQzvJk8IsWX9SQavN2
bfKILRGJ0pheAmSz97yyGO0sDyTcgoeZYhyWhP0BGmJie8bCgdp2pIKmiB4IJQBR
3r/IrAuQCTH7dK8iefAVcqIQCwZZeNqtRK9hxFrhTFkoMB/wwwk7JP1ENPzVtYCE
ichNvQhNHJzZ7eZ25PeL3FwBp3VMHqXoBcfZaOYx7sR7C0LBXU/QbUc1H8iX/ll9
iIjXJZDKj78I9fSwAU4p1xl7xqp47l2lViINPBhrgHxaTOxTTH/j3Q8z0BnmwDFS
E1S9jakSdXyTUHj4og+3vhIu171LH5003kPdLGhrityRJySjmXXT7yygDsKqeoVo
i5aB49y/4jX2GyVO0HYVDUlXInOajYyLvVpme2P5MqHlkd9IBdMpgIIXwxU1O1BE
ywvP/VC4ossIt5UOImk8ZuNFOq2WrSqmjM7aftoY10yz28X8NDPddErknlL8jtMA
eTs5dA5pF/Zfo4ucgRoHWuNUIzZgy5X8rk7cwwnjgNeewrKDruehA7PrN9DvFgDV
Ei5cAc8OqAwG50HwK97mq3PGuv84tcWhBs4KR6f6Bj6+noMv6TQrxUOUnqyFfckA
iFpXllUmEG4gx8yyKcXVUtjJiQiy0k736rVGCuxzEypPUwoIfW4FnhjLtp2mS4Wk
szeus03E7KemLRX3nBa89MG7AxyERlEA8Fh8Il9NpGdlYZs04n575SOyuPmJ945s
11Of+K8FavoDwauX9qZJJp97CFg4etBEt20JGApc668mcG0W+duJ1vFjAggs3RR/
UGTKFJaOW2ACB9xmRZHOQpHI19/7VyDLmTQRIQKltdv5ToukUQo8cOyRS0UwNtyS
JgblgAfo0AeHaP3miOVZQ3DZ/KsTaNvdpU3R76QqGgmjkukfNqPo7YuGMKb7+Rj+
3L9DznphFxzprYm1uuzX5pHEaGa6GQ/ihU6CLYEOxbHJXNbFkRa7YUxM9ezD8wpB
dAne3tyHCdhA9b8Tz1bqwAYMFKz9j63IhxotDNfxQVd9z2UFIBB9F4qn/UfiG1P0
qE4jN0SyW2KjisRKpJpQXWzQO2uNx5+E3iUmxvMYeD9t6zYfNTu9ham4378LOyO8
X0MbCaz8eks3lwgOkQSrogfYmuP8L85FhEQLf1BeUgBcTwoJ6awN4JY6yuGlKQDo
Mz1sUCL8Di7eBNkrNr2MNWkQO3OVFoN7lINfeZsw919B78VJxbusmwdecD8wUaMt
3TYU9KkYa4YBXgY2VlZnLJzWYl+zAXnIzZ3Dk9BNf8XTWvqlfb83bRgzekSpbZSb
1aSQu0DqaOY1dmUNNw84ogb8oBTELMITWj4KV9PpQsPWy2YxSrkx6STJ8uuO4Rjn
HhLaaRn8LP6Dnc3OhS6eXEV6nTEgE+D4BvqG809JtUOtb0MWd/GGZia/N1ckS6ZM
+PQdQ7OTr2MCpGJGgYrmOFOHvR1EVwrt0DHSqLG9M7u6NLAxipOhnJa/c8J3re29
16FiOK9/p9nEcmvEAcYkFGVYLvotBhNRIxDaV/0vZuND/n9ixggAwEabRQ2dJ1hO
YSETa/ZHhRda/9xTja7gtbH60oFIsS+2GFltyFO7B4ni0YWdZXSsSxb8DtGyYriy
8a2dVS6vGX5qLPiSnjcaf6X0Y7sZ6y1XrGzV3AYvUitnTxqJDmrn94TNDfjigUZg
G0/4UFVYPN2wbfXYk3y9s+LMYUaYmo9K8uorg9ojbo6ivvUigf1Kzu4ogW5KWYKB
aGOHDtavyoMutSRoeCEfMgzMvQB8mBy9q704IJo1UMOqP35IUj6D4Mgd46LZ/6t7
5Fc354qxegdcfDO65grN3rtBjCrZ9rNqOj1OROwMi1fuE1t8H+e5kACmqOZL6kpx
qwGKzi51rzXSnIs13c9y8U2SVOVZdKyWcVC+PJLoc2MHGKZNZqhYGlmrZDFIwtZ/
5s0GwOPfKn0Mn+dwPVccJz5RbUBO8Xz7GxHobvJAI1M1jB7/LlEOFDdfdBsij3Uc
GiNaQYsGxHnEVqkDKLlC8jyscBOPeQy7X1k6GONQxHWPE+BIl2ONGLgC21uXDZ6U
9U7BytrKla8kgUpf9DU43zInjzXv5H62b+EAEwDil/3eV40McPuWpRb3/Ip+mvJZ
2qlaIrhQdiHz5YOKVq3ACVxOEPJmpHnUyHemPZRbhOISqBCmYYVhQNQjwHMVHHjj
DOkb8TbGLncreVXL3N5GAuWh6aZBDUjs/DKD8KmDBP5zrp3gxjRzihHJt9WutX0s
HrXiHwYWAJaMGv8cAlHvfo8acfYquUx+n27co5GEbewbuXZSKl72WuHsKuTwUVpv
52qymb5Xrq72T4OVR0Hi1AFkx4COi9M/l1lK1qrLMzhmsWKGfLRai0fVsOCmXMRD
Mv63LwElQYzaRpDNzCWEdGHwZ+U3zksy+q51J91mbae4JM/kXNIHapj5VR6wbWUS
LKMUKvM81SRV3eSzZmLEqOZzGtB3ZZXBeB4w3WSB7L3siaE3gPmFWeT8B5sqAIAj
esYxMHx24Zvf33hBwOWeaplo/S6PX/Z5YjtdnKLsohRTRs5yt9xpXeHyKRipgzE2
/SOkrIOrBWEomc8vcIucn7TU0yUZjix03noyBMxGJ2KVsx9YcHzTytUCovwk1KWd
AYPvzWRlTBq+aylNuvB8iiVDXSplWAJCWOGMHhaY7PkaYHsYkQVjdl1J1Gn+UPkt
HESUyUX25gTcARw3iIQ/GbElEwuPsMzR+mXIQfLMy6c/RebX3ESnYRPUaSVDASc+
haT9YEvb0SYKE9/2VZVjM++l1GLlHwIbZSBNNet4POx9WlzIelS/8Q2mjVa5SWym
mGSZTfraW5X39BeutbKKJ7kanOwx8dwl9YsoQgchFiTls1ubcBWPpaAgIQ4kjNG9
/jIhyyxeCGnxYR/ITASouE+cQmEFJ0Vk1WYn+ipzSrsjmfaqZnrKVAptjdmppaok
ITwWmERd0ZPfXZPdANdalGh1pZT1Y8hY295bI0XhaukO1wRmIHi9gBZaiQFkCLBT
8ojRDz0OvHOs/Iinai4ZJAKjViF7R6Zb9SyNJpoU3Fz8UYIdpLLc8takJV1wRYq3
TgpepnV5Es/DHM4j52uAPxO87MEo1au79Y95xYTDyynJrSkBRasXhMakMg+PqDi8
pEolcyncKmOE+k6IpaLPyqHxg8TeP4yhCLV5hoBHj1RKHXSTfvtOIkXd1XMqLy60
3D+WEyrA1AWtRM0ngA4NJJ3C/Suo2bjxGsD0cmFN4qVSOjpgjSq6R2vDJ+e4SdfU
YMO1G8ZzU8eCsHzealtn2rfvy6LrWQTr87tvD9JoriRwEFrkGMecEqRLag09IDM+
Rh8ixfUu9syYaQZQDxnnhsw2ekr2C1S7+Ce/u944S4oDDcAbbD85sU2bB3l1T3gb
sPgNBKCR381lmFUYWyWUCwtN2eKp4qQqnKa1e0NWZYgoayOvLooBQBp3OR95Z77Q
9pagTyZiC7XJ6Muo/eXUEw==
`pragma protect end_protected

`endif // `ifndef _VSL_MSBE_SV_


