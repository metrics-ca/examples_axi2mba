//----------------------------------------------------------------------
/**
 * @file xvip_axi_lock_scen.sv
 * @brief Defines XVIP AXI lock access scenario class.
 *
 * This file contains the following XVIP AXI lock access scenario related
 * classes.
 * - XVIP AXI lock access scenario class
 * - XVIP AXI scenario election class
 * - XVIP AXI lock access scenario class for multi-stream scenario
 */
/*
 * Copyright (C) 2007-2009 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _XVIP_AXI_LOCK_SCEN_SV_
`define _XVIP_AXI_LOCK_SCEN_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
bF9VTSNvAr7tshvw0FGLTuRIhwGDrjOVamTKq5EfQ89AGf2oA2oBmQqa3JM0y2eo
9m2K5xt3vVnGogvxQByNWOiwVXKyauL4NoqfCOizVg4iz/LdC1CLb09aDswaYnZ+
MhpvIE6RK+Bhz2fJOzCwqoHrOrXBat8dWyH5zVwtF10BVByeSC5V2lm9kk0SlX7a
PWIa185qbcQNiCEatAWnzU4N43tt0Noj6EIZGtXn7PcrJRH0dD6Nb8BpPrfQ2yNg
SqDR2iumRv/t6jChrDIKAikm5oIZxtDdX/aQZOuz9Y7G51iNQJ8w2XMZUGON9FaQ
jqbXq/cn7K+egue69iTYzA==
`pragma protect data_block
j54RHIrA/IPZ/QBH2xA9HJe29QJhuA8FTQF6LTSwJ69QKTunuGZSwhxXn+dbq2kx
mUEn5EzcHxIxSzFmJyRXEQ2uQwUf2r79tjnBv7CUmUzDcAKDQGZ5rz9YEFSlTb3s
LUNQ+aZm5U93TpIOz7CWqdOK7B4eXNVV7ieZwBoEL+KF6JelI/tjQeZ3L+8wxQy0
7bA+8XS08rCkpqNIj0rGo2elGBx+RbqBAkHHVSCpBaE8GQj0E2ePNzxPiwWiqT5J
6yDmHxQI7YXN7gvo/QlSmP8maC3FeIsXqtIxvngZV1Twf8jC0t2UHomJlvsv9AWg
aDGbVl+z0UVjJqbHTRCEZV7ssGRBApHYPxfD/vFGr7mM+KjpvW+mVIcqj5ZTK7rC
zqvp6pEICfmhWtkXziHszQX6DI+1MNYxX0jpxsdwqdiUyENd1FAI9s2tzoL4PCj2
6hSRHe5VZQAQouqDoZTQ/lvApFQjOciQK5URGtPpXcXj3pM41ThS1ZOVVdbJ8PmI
dubZdd6XkEO4N6IVMO6koNpNqb7Qo05q7DKjiUKyDKWmvqGDdRnAZIT8p59DDDYe
PeL0STkeWqY9k0PFSZbDngD2Cp9ehX9sgETZii1nTQSKysxwAWMe5+0c7Qoh9dJC
r39nm8tvqHOgr5ZMZ+QPqwF8YyU+hXbuhRrSaeK1bv30A/jV8MhSgvmsFsTwE25N
YquzGCA8pckSY/dm9n1wqwtjqpGRmT7A/w1n6WEdZqx3v2X316ow4aQo2CDSQlbY
Bf+KcD8wOUkR7OofH08UPGXRTvwYXQmGTRu1N0zHsh9LEUZ973/ULsFZJfc5Uuf0
5lDQfzc8IeNGZ5OlpyZjraO+7uSODDIUTFZ/XTFmqNZqBfZrFeyjhJ+cXk1hqTUq
unB7kZA1u0N80p13NFUeFNssNyf4LzyrkuaWzCbGiCC0onn+KtHbuClBWtPRbRFD
YIJEf7b8RX5f6HXc3/rSw0NptY9W25p9YkWTMUf8p0nG6HVJbc6+/CTT10upXlEA
1BBbIVF2z3Kf3lK99IY72zHY2L4jKhlciz3EaIOmszdTB0RzqyN/q8C77QIR0SSJ
4rMUeYuQyl/eBykEGD8QHZlRhYLUFo1cxWCxTyx7OBM3T1Sol096eYFLxuYPBQ+t
ouPgo9PeJB1Iel/Msjcef4KVpJapnLexWoYjrhO23FImpiGVvyzu53tn7wdc/U9e
T1YUPEypMM4nszJVVsSAfivkxiFBdPGBwwdyWlKtNleL0darp2vGUWifmgxW7rIb
Bd+cJlS5K03n2t9JlumAlqyb9kJXJHs+k3UoN6XYVzDn83YviNRDBaQE34DThWco
Tk2/J1F7sRM/hATnFOSpLxmcVnRoWyQyUToRR4C1CHRvRNVwqw/ZPStdEyrzOUUG
KjbMTiBAUTrEW3Ces+6ah5dOmN3eGdweag8KmTJ3nu2OMWp1Rfhxa5SZnsTwIqi3
787rxB3YjFtfy8F287UFEYBlKrHtDjkThQUNXbO9+SKk6tL+JC70Zrix1NwnZncf
NGTD8p/RkSTlUGSop/Hzf1u7e8ePS4Maw11KJzpQO5RU2Ssm4RZJXpOqgecDIG3i
l2dAXa7k+3TWtNxbTX/iemRYRyYQ3yYmGJvg5/t/DC5X9rBWojIUONq+Ba/cuA/Q
k9dbIAVvhWDCkvZgrBlTQ5Boxw8NQFC8xAu5NcTuyqQ1zfkka0UP/wRpLsmcvsHu
L67mrP0lQAFGQ5VKWz95e0vl9qrUjMajrDpk55V9WM6wjst1NSqZGgQKwFr7ttNv
N1P/MxPRHAIFcx4Vcnki3K2KXK0wR8foQic2vko5jWjO985Jt9E5imK/ex/LPXdO
1NVTq9cKNf5C6/CfgJwtVF9ZeirszbUeWjoTrHf2qn693lf8YUloOXxszDTJxSlJ
NToLsvd7RpxK4fI7lUB3VA8ppWKBpwtXh3ufiefKNsLw3vPF/2n0LxFLhT77fFEj
EkdQFR/Oper/MIBwZBxziP+p44VwgE+ff+4SYeYFkTblZw5FvUKFPJUELzLdz+wD
aEtS02i3lDXXM362rKDo/JIs5H6woXgbfFmS/2QwLc0qAJf0b3GPY9Xfg3E9G9Is
lGCRcINIrC7+mT6ultRgYCpPrgDxxrwuVbPVyvoWnbnJwVFR1qO/KKh/mHG8EJvt
ZvxupWu8Q1pVvO+POajTzvEafafcwtVHhNGvi6viSeE3DL1M20RS9xnS/Xo7Fvjd
8zMKRjsru6fsJ4r2Biz0nyFCVuaiKtl8bRDq/M5koyVrl3Wk3L3ZQnjs8Ttc3wRH
7W+JxeExhawse9qxwI1OyybiVBF242Ea9smIV+YIYrtI0ypcJ21Q+JEiPkRMwdNS
/hCZXtyxGYR6fT/sNr9CNYA8oKgpJ78sFyIzl51o+Cx3PU27w6umNN2+BCcEsw7K
zZWxZv1SuEjSflemRB5AbroxBRCTZYa4utPSnsP/JHtJd5tg04AsmCXsb+P6X9lP
McXAR+cPooZEDi0rbon3EvACMtMNiY/bcB0GILOss0nPLOTqy7+kFvus9m+ufnEY
u6wfyl8t1V/z7ScxYIxfUQnmw7RQJi5+2nJDBj9vQWlrrZyStKmc/bNepfqN2OZf
zUREuK7KOCfFX1Q63L9//tyjvzm5cBkWR2RdtKOHH8DigSOpg2BITjB5DT9+s6EQ
28wztUWJr1lQtYL0ssSC51n4hyc5XeuDVSaZQ3FnDymyZann7eYovphhnoXc10nL
T4tOud/iKaCmQNaVcbhWP9w/paCvn2u8kQrUia7flaVz7JXPGQ2sX8QAjYNKeyrb
BPHfvH9+8alcMPgNxG4FUNy8tfPldh/+huzWQNsryXJm4yzV8EqZjYcG56pbNJfn
H8/73txmx7ImohoHn5QUr3oz0qas5DDpmdFgarS9XTnE6h68bfF9WwsayhUWEyN9
lSmYCJsbtDnY42+mLIFX8+fFn2E4GE9K8/ZLi05VvvwwmKCQtAulzQF54yjpU7mv
BQF6ubJP/G2dxHNiRi0CHZ+wMmn9IFXF7NHnY7B/LztUnRrIA36oxCAOR0J39Aws
fo9VRGPIFz2MwsIsU7zOXNqqhNg6qBMe1vbiu+Mt4Wioj8OJtGYsMk7kKlgXctr3
o9AG6QemTujut1ndZ9gHFeaQTuw+msR5XxazksiFw/QroGrussodbMRh4Fc1RdvV
PF15tvNRShHfmxjFGDeHqYzHAL4/LH0JR7pVP4/rwaiDvXRc8VhFuFSuIlR6VV0S
YdzCo8vimTWFg/HC+V14B8HWai9qYI56dsJ4CuvyRptiVyy3hExG89acUv9/EOUP
In5Y7KMhMZcmi5zh2JDqqSw+nXI92ZnhRfUAGzt6zdkxY/UARFtWr3cdTZFRY9aU
hZmPeWIrxUwxjHF1loSg4sLQ8dj/szoXY7H14UauSLftRG+U4tHGsgaS10hEn71n
Kfve1x1kauMMvTVae9lkp3ZlIheJIsHQXwfvJSub88+vJoKW/Tb/G+Ofg0leFWgW
6oBYz3pXchAfEUwPuODtEhHki4UkGptHeRm7Ha3pA+LHmzEeaG5wMmpqwj/QGClK
qLcg2Pi02jKH3B3KH5I2JTPiUCVaqfivdUsF49+FM6VM3HqbrttlcqMvTJOxLtWt
MoslyiRpMZ+/wh9RHwPs31BV/v9XFlYC66dlJsGyf0qGbEBeTisvYzxovTDeBWa8
lcwMEW2ziFCZMexFWFhv9WGbUqq718yCyUqI7GJpaHmYywfE0s46RIThjV0Kbwu4
PVipEnXcQnAsoJW6LTsikwIDyyhoQPOsGnSGYfVB02WaFs3p/hh6Isqun4TAojfC
WxwIKBLPs35JrXNt+Vk/6Md4H3Hx0kfQaK++dwLVWbqaMxKc1eq1DM7x/Qh6Abxh
xPUGzhRzyI0PGomsj7JnYhm5urYnBF1SNvvkCloUqcsCuyP7IyFdiwIinXbSNW3D
ihJP7/ZQzZLDbKLM1qFDHFkz5I2xZFMeXbErKgFlZ93OzPTMGn0bP4k8J67ME4OE
OauIw2/OgmR668qjz2NYJ8nlIBg75ypJFDrKN2OyAZUkZ5J040DfVJOZp/Y1LsZB
VUy6gnJPpegU/V8HA1XUKnNzHI2VwT5ZqGtS8MPJMkwjnKhLh+pnhs1k54xR6Qdz
mtyXUJzPT/+2aIIB2/6tlPiVI8nY00R4m2AEe6l0Wb8qJsZouVCLhfihPB7JySLV
BNbJLsu4cEAdxlFtapnfo1QqCBHBNg0hc0jwUpqWWg/owy02JbxOvFk1hwWQ483f
p2RFZn5OJFiL4eMU3Q1Tw4NAgAjOUiJzLpP45x8OW4L2z1zOboTyXobl9c+J88L5
KBOQFD3/ltOuKSqOVAVptSEsHJ1YXGBNUyXxbfGvlo3Ig/6ZOGY1WQd3ORrbOuMo
tFbmZBcjfNgqXxwNeaH0c5MDe79Tjy/6Z42DYgBXiNnmByL2cS7XjjWt5RiPdGaG
InDE4Aol9mWawTZY14Hv02uArCSU9vt3OM+JZKX+9BiGLRDOD9YwJEftJO86EKHl
+MeSKKyUsv1Alu6xHRwDXxLPis7xGjhcBxkiBUMqwhb5oVwnBtIWvpUQDr8GGQd3
4n0NP6AxexH65PdXFq/wSvICgObzYl2C34AJh1/ZZOnq6JrNaaAHkifgtk0Cf4rU
Fr2Q6eRH341aK9cI+KTU1FZmiioFY7vvfI+gIlSdDcpp760sY7rxy/X8/r8mWLBI
9GEhpj8PbHSyIZMegjWU/nMOmGOhopipNRj+8hAyAjUfysDMAK9jEFS2+D9iFlFu
YIvUingj9zbdCvOX1wfTKY9FIEJ9Y5kW7NXxBnpQQH1+CRVG5uwVyU0ZNCuDAEeG
ZkUSSSOMWvO8OR2ujM1Frx/vrqbUW0fUqvY4pSngAwuB3ShkYBLpOOhlf8OH/y72
HYtNu4YulMgWninCqh+lEqCjuq+K2lnMZ9k4yGSFuJBEJY5q/5/RuAwVBzac21ox
Acpky2e9JIY7+TQKgl8URWwEpXjYJESe5aUK51+BqDLqpfomXhyD38rdAw146r9A
pq4pbiIgYrRb/YLluoifSfPjZdC/fuB9jS7V1K3EZpZRUqk4Jc74QujaSHpcTJNt
uKaT/Dpahsh19QExtfXpAQK6O6QMknDO39Uop+wkbH1yBhCUlDbhM22F05MBrRom
shyYSIp00Q9blWmxH0AXPMVuWvGmPaBQovqLwL/p7eYxO1j4ONlNX1iW9a6z/5C8
UfaMPXK76o82ekznp8E6Vu5zcfiLHGXHjzlc9++8gnomc3yyPIW3o9Zskhmg/vmn
ZsAVDkImteVSLuD8qqBsjv2shApqGiNLpsvuGw4RsK2yZ1s9V90MeBzgErj9JiWE
cQcSE6Oxt0bCnkJ44Z9xQx4sNPN2rkp81eW6Wa7QLgDZKAoUPHUPH6++Me9XLFk5
dXfdjp7q8qBSo+rqqqr8gqWdARG8YB+k8aglV4BvZWtmAOoGU3QYH/B54gUA45Sv
Cjn9ocSZST1y+3d2RPgWIpIyztFy0KA74iswnTapUL9r8kygkyhinZ8/b+fyDVGF
krxtxC/uG+wq7gbG6eLcrJPbwhioEc+DceKoQM0vbvGDRDtHECf9dSNh0xVpJlum
CjylLAUryTmYa1A7/MqawLKoXbhxI3k+AnzWdu+QlHWkFafgCPCqYw2f5UV+FJJ/
VhCCBgNgwFMSPA+vEiG8vQxNG6KCo48L2qsuC7f1FhzRbguBti8N7+1Dfx0o8fI1
N22jK+n0Gg0plr5G7YGK1dshwvC86zfhPMzdmL6pnWUAexQo9MaDoD0gATR7fmZe
KX3e1S2EB4dLrPm4vcyH6I0vti56Gw1xJ9HFaSsh6By2TyQs47HC888Ch2oeMoki
M5RLaHgiSgWmW0q+2xjAK0jCmTwxWxoBFrJTSKJCFe2FIHpI2TOJGUdV3inWlEVV
tt28coxTUQu8QkJwcVpDtWPZKJHwKF2ihUlmIgROvGhyq4bx+QCDTVHVWXb0l9b6
T8VRpBt5nNhtxxb/JlLvrDZJzZhklc0sDyq/nopDKnxLfJ7OxqyDpUqYh7+6ENvw
mNEoGt36ZkKaW/wdfECYRe+qHkw/Nw4PfEbSUCB+44MKX7vZPhdwn7/eT1nDz2k4
7154otgdaxjAXs2YflJ5Ttq+6xezmHSFWWz7IIZY0Z5+zYhvfU1IP9Z/M6SxqooU
X5rs0fWOTxF1fcjyyOMI2QeOB+qmdEvoXCYzgAAceGZUDxAoIGcd6Ndlse/3R6r5
+X74GxK1o2pTPOKEIOiLgC+gc6mzYHUEyenodUx6URW95nkmCdFolDDEQicRNngj
oaKCjh5j4i1hfOvVImdpbhno0yM4AG3yj/2veMpxoNCGLl7dK6ywianrmc9oVZFD
V5W9WDBCMETm6l0jyRq5YvdygNj/38nfTxu+3S4hwEazygQYgMhRgD7G6660wS4a
WBBVZhLlRNNDHq8Dp1efkL09PUzcrTMvkDKQj6IL49AylsSsSS7XNPHpCgcl8mFY
GaiSojqV3ZePMoHmSU/fetCV56sJwe6efg1xGZKXTksMjrXHob47Ln/AtdwxCsbq
YNYfRSPmDNyjX5OtJNxaCLF0xloOqTOqVW7Pzh1ljtIMWkrklZkrKy7mIWv5Kb5s
jVBYSbDwTHd8CwD4/qKI2XH7H3whiqA/jTHz01V6DInS8wglKxVDGHhyOIcVb/fo
YDkFhZ8LPCKInnZECCnpB4dQ2Eg9zrqO3d4DHWC+XosTk1Skf/izjn+8x3JsizBl
f0kF3yxFQep7Jzwyp8E+yC9j4timAc+3QFoY8NazXCMBko1FNBLUnGxNiobuILMl
zXncwnqfzw0mhXemGOGEMhrkxvcsPIKBr3/eheCqwCHg29SXnzIsUIiqDYJjSdIS
SMF3KwqjufUu3dCbV6f3YOPWVvds8FknEFKO5CmAXHMJW6FFpfybDo/O/b/ZqbOY
bK8qCmOP/zczNSOgIoVcxcmu3U7DwfqDVMcoublUFBuTHhjwtZnQzX+HWyE9tJRX
Q6VHarjUaXcMMZxKKCeQEbum3YsrrtLaxT8Wav9nwgnxOzoyMXEBtX/xcCBn448+
IxcjOiGS87RsMCAZWOGKw0Vm9f7Nv3CH2+b0kyVkiTT2q9RuVALAf0sQCD0aqynU
cIXke573Xq7kedwL67q4tz/qXvL3rV7Y5Rr+EWf2oTDPwFHlHQnf0FmQOrUcdEqW
i4sh6WZChLglGYlScAOJ6z0bWUMtDyoh3N80ZTSq443jA3iRPGDHBvHXH7trBkXB
sRKcOtr+v9zgOk3JhWTuVRuMz21QS8+6mSn4bIQUFYabZPnvBnGTuxi+GAUt+1Ip
YCsVQ8ec33UzCwFatdjApyFuR8twsgvn5vDp/AsgyFCFRIRN8vKayUTJfeD87Zjd
q4a2VJQ4z0qIf+DZHC2+yrhkVsVqAZ2dWCMnmvmlEq+OQLJ0i6QsEsAO+bs262bp
7vJ8EIoIkvbsSjmgen3z+PMIO7D/kf2wYeUMK3BxkJr+ayIqmnMF+PdFk29HP9ic
5utlNBzp5Mg9L/EjN5BKxWJqORzgigqXrXtLLMLmoN8mLiHRQmXarzr7Gp1/wvk2
UDV7uW+5RgLpqhSO90zt0DoM9dYjlmyMFdcU2V2CW4Wpun/GfZEbOtUKpSXKyOZB
wB6L+ZdEXjrVL/M9iuCaofSlU7xf+peJljXaq3q0Z/lhOoLzKqOGEVrT58Hbl1+4
nKTH9EsKtBgKphVALbhxyxIvJakvhsQGQAEEt5v/6Wki4oMlrF54XhSPPOGho7d6
6j/N/4eXFZJUwBel1/DMIpNdKjvgWKFTk9y4muGQwc+j5eGoJCWGMAUPb6GfrOO9
IM9LmjLKPnCK4D4DrBAY4STMf2Ay1PmEpuVMf5a6maPBs1GEGqkH73k5bDcAZnoE
DpEGLSvgh49Y9fXp8Zed7ESeniqfORn260r7wDgXHK4A9hzaLFw4Wa1jAjV2SPdp
mNlSdxbLQS2imBkgyfio5WZ+Ivj0t0KSR8XROKvllnVOtq1S1APxnRGw/tlk0tQc
1fOHq9bBZDc6PlWeb+oFykMxylj24mILLcp5Erqh54SQ+4fecwOLUlopk3fw4V1p
S912obEvII17Fyo5Nomj5JxiwzH0oW3tzFD37n4aT9SLA6JEQRHEMqOiW5gmJN59
ED422FeX5aPDqOagzIUL6NTZgOCluNDIkf2idkNMhAjrA9ptkrWU66+mdMOPWkS4
8Bu0ThN6jBt71Mgn4T8b3ObVA5TQEoNcUo7Pyu8hbWhW1UVQE9StwTqRD14geYRW
5DIJEmNFuxFtGlu2FNw25pSRWh7cMdjZnXBM5REExsGOiBTm4B9Y78TH4B8/lfH0
WtCEtOdZy3p6rGME5NiBhsEhHvca3zaV1p0uC37c8iVFKemoW2hKmIqB0LN3XN2p
LwDkhPAUECpj2f9TGG+gZEoYvwU4vRTuUdljajqf65Db/ZNHs6u97vKjDeMTTRAF
nR9zI7XguPtDjmyLKPPMh4ayYlmfuCVyrMp2GyRHkpEyx6WWFlppNBikrMJ8cU9h
IIKpdVNBeC3khcTXnT57+HXzYB91tUGsJPStY9J25A0EgL2supDCFOeyVsjK9k1j
virzuD5EVJXeLK6/kGYvqGTj1xP8ARQRtupYQsIUaIHbYZYaasg96ie3avMnDOYX
DrAE8CP3IdpxzXjyS0g5S1d4Wan5mVxw2pGfEKiXngaumr/xDMd2Oglrf662wFwV
Lu6OqjjGoImpI4rQRb1FxYIMbqS6+ZXuSFKx5g2WgQCmrFuHsoQ4eZ5RLCMGAvlX
9rnTzaRftZgAjYDLWgyPvA63+QHSHliT5qI4OFdxXNOXmE59Wkyu05+827ulPXF3
8dqxuJ52VNhBh/vsAZBBfYkcgbMMYEMJYj09PF9F44euWvT0QsDrSSP1bhcOT3tE
X+ogGHjhBlbr6rmkLDLs5CGZ/SWrZwX9H044hwjCzWV1+t0Wgm1cCDCx/o/x9nPu
x0zba4JgVaUIZxY9cB49t3wmWOhlbW4TWUY6qrP+c/lvkvljyIhQFcjR6xdbhLdK
aHxZ9/NxSd2WZJIo9ODJw66x82N6K9wCT2GOvvBfZZVoOy4InP35RC808h0cz46Z
x8ajkDR5UeR8WN3EPEimEQn5wntlXxDnTlCd97p/QaS+zhQii1mGMceGbR3yYF67
1+onFjbjB+NrdFc4AvT0vvSidkO5ySqgp0Rj0fJwOFbxO4u7oWfKcTpBr8IA9XX/
wJlflC93p9GC46Yl9sWkBRxFbpeKyCoLge9TmktCZdKdunEsYtA1bc4onshddwS3
lZ8fJrKx87p48WnHvKtxSIbGY7pYXUmvUB69IM62lmCpdfetKgtjsI1FGVSaGdkR
+vY3eN+N3dcVxfHP6YrT6B0kEoqKKYEpbZy6WC493X5nCfBJLCrph7KMXeQgmZKK
YkDxloRsddpmYOpB/qhU472YKeKBhom7L+/7pOPMLkiRADxvQxaDohfdF1yfWeH0
Y5JT3G4Yklj7jS3lOC3hhOImRiKlHbZxRceicT1yg+zUJZTbOMV+YSUxbFHcHxSa
R8KwqL/yJ9KdVK6OT41yF56Yuxl77+uRu2wJjnnlD/AINTLSf4yifsQNzIAD6RuB
Q+WIfe7gjg80eVsLJFZ4v+IahE6dLour8OPBES6D9uvuHpBTBk5O0KtEwWWeBfWA
IG2PF6I862T0dgIUWScHVfsAAqVX4gqI1QUl+UZR+bgkITBZgAfgNgNy0r4agYo6
Aa80CmYba70Qwh7K3/76fr1harQ8E47WBhkTnuue3nnijnRKKD3zwIGRmp1SrKIq
HLllO4QzCyLk2m7QadlY3FMffOSpDLSHNy6B6v9uVGP+Sxca+8UYhDHevBfl3An1
JJ/WdqlOuAY1Hkfcpr0HqFAaYc33p7vyZx0E/rB9iqz5shXXXORXclYJbApl5vwx
6zZUpkYgaQjkLTzUzevG5gU7ymJNf+ZHvbr3nuOUmXt4V6pekU3SH8DtSJTAjPfy
+RXj8af1yGCgqkwQkHEAW1lZpeKuWqVE1Aave7Vno8yC5oYLRnwNPJmAeBVKY2UN
U413XDDqrsNm6KAGZL5pQIgjFTjwBUagj0Zq4g3z5mPoo3Fu82UZqllqanu0dcXB
0Frgk3paS1SIH176EweL8n5O0BLy+YymgNmTEBezpr6qTchf5Goc8rp/0Yq7mwJc
/Ewv/TmFkvLQtuuzs+JePyQFtvcTNQOGEFdEHsWxzM+IpDwWskAW7IcgdEmE1kNR
yLCZXHXzlbC+UhKoHfOQbGTaoShbk8gC/B9KJPMjcyUHCZ+jBhG/NIPnQSH/hs7M
UChbUwt98DzdnfReWkGGlM1KzY2fVlwoZD0k2PD/gi2cjyeDrt7EytEoW1H/s1Uu
nuLM9kKFA+ZmTQehMaimz9lC3J1nQqXCD+AotbSRRAuIIrWVpCvyS2WeGLH4apwe
k2dPAnw8U0uw0cGT/96+Yv8VRcq31LOj8/0lLR4esWGo24JjsaZjRChlaHka/eIc
yKAvuDVhOOg0tPyNHGdUhdQ2f+KVcgCWj4ecckDpx0S2SJYapGgiRUKfeMn7NzBZ
jc9RJBqChNcJyhaBozrH9/hTryYou+x/3x6I/Zdbqcjhkt6laUtS8wZf0NVWzqe0
FrOjEgXi740hxU04tBcau3tSEH1OUDbvvNJ0HLy3TWTWbu07rWu9hg4rnSzpNgPM
ScGPjlGEmchuUMTrHz8w3ogXT7UhLL5//8hltad6T8zGy9OyuwvJLpg+KjrLUqzB
mRPDMfHIBCxE3sfG21hP5ZsbZUYvepuf0dRjR1sPSUDdmVZzw15rJwimy7RuX/0y
2FkJh1krmKesWi4PyAorwUo+tp4S4qLK6ramjgwHvi/Se09RRq+svY237EOjFtud
Rk1jlUxwdN+WV7xBHpOvQJ+O1R8OxwvT39mCdtJr0dM4d8c87BdZKmu3eLj7Mn+p
cHURakiwKHvrd3oU3/55Bd24FI6kHAMoSSL8SlQcJW1GdC+NtsbGb6j9s/FdbuUx
gV/nkCetFT4X96fKqn0Xz2gHbdPJWwxeAncOJg34DKH0KE1G+mKcNh9zqRQFU9F4
yEFcS8xb85k2+BHq17fAfqvCXpvv2W7w+YSCWn3ljvJeiKWv2fGBkRoCGZBR0Td/
6VE7RjDhP1+kA2xG8h3BMjf1ptFldXHq8KWGoYZVAsY71q2UVZsoDg03MMAX282z
yczhxoR3nzJbs0TWzJISzgy9YrS/IRfEOv8Q7UrPofrSDFTDoWQqAUaWHvgAL/bd
d7vI4ONrX7KRcJclzbzd9QA8qiMd/zlWei0uX5aD7jg6O3wcJ+yP+mLZVwbDwg5i
BZvy/XUwC9JOAxj9Ehnnu2lbHgNCcJOfdxcHM9rZ3/2yDjqGjAuskt3ta3NkYNuE
0D3WQp00+yH2Fim21VRuyg2o3xozTyeQ0EPsvpwK7HP38Rekis5Ck1sTjq5kkSHt
PNl8xZk80dm+RtqWv8jlm7ISojybC763l53GruufE9Ij1aVq859LyVgxgUvntfWZ
oJ3E8rri8ca+eZ2cAvRFaKHQNdXP0vj/hgAV9OEvUSxpInTUySMEsnQ/+RNx2DNv
2jThIS4rGhZR21sejN9rhiR1eGRMyY4pCcXM6nNNkJmox2A4d0RtqlF4KhiNojxZ
dXdf4c1rnRlBIg3wfVYc1wFNwbf1kh7e6LjsiYTCMhjcSYnq5dlyUA12rOXFoQM3
3yzxn+w6GFuw/daeIEtu1u9dKXRDLV872rPKFM61U/ZE5+R/wdWnG60kW80bXszV
1F1ljNpT7IcAy9i2W+s4cXljCiB3T0JibjLa0TwoQuYMf1RRY8qUWKPpGzpB+9mx
k6DFqK0exkMWspkv6WsBMAm752SRDHMv985b4c7e4L7Q1arX/0qsdXHD8eqPpaSx
EPxIk7QAuHFbMbFcub9wOUIZo8Fay0V2E4zxFQMtXaFZ7ch68tn7oGa83+K6Gq5L
x9JjdH+q7qpQfwhcoeXtN1V8pM5YhtBdg4XQwRofQMc9uQpyxR7PWdA8gmobcIXM
l+nq1eCMMW3JViIuL5LSkfWJSeRDHXS8B6E2f6mqNu85A8W2/h7rAhNB6ZA8DXrn
Z1eID9T1bMtsD06G17KF12MR0GUALCttBUH7bOv1XnbGqxZVb6nGFe+VNcg5bCeu
jQsRE4xg1IZLkFoQf2l7ExV86RSnnpBr2znnoH8FSx/eGKn+DTVcYDOoAOgwdGWT
+x+0Px27cvYyUPnlEn6ZgJvFJSxeN/DgUaq/VKCptJ6anahm19p2l0RA6pP09w6P
doPkxbIbEri7mOuIFYDAGNmMq3WTrdDBrpTqGWxnfjt+VCwzNtwhDmaM9WJJGHtR
b0cxfNtCTwiD1V1tqesJWnngroN80c/o6XlvSUaTESfsiB8baPVV0a51yTgH6JJe
qbmJhRFBdjmq4d5EbOvuPO//J1kivoQ+zRoJqkUu3CLID/sZHAuufLosUHGhNJ9H
0CxmVECKPlJT3bHpYMVLRO6jQwPWjEgNgEYW82kEfVqRQ2jYf7F1/zWf38kQkECp
64/5Jt/TMEyUautgHsKBGsEX+7WLgD9/HMc2y4deNDIlfzjR2sBV3uywshYM1loe
vUEpTNRS2F37h60FuLZrXcQkTcxGQ0eVC95uF9AjC2GIE8M30zms6pZEXec9ADrF
i/mvELhox46oEzR9x6G3hwroaSNvA5ao6E4HSbo1CzQ3BT0GT+85pKDs2DsG83pG
O5eDDVOlWcMlrRv/zCeiicdSz7iJyCQTbVJ+IrrUwJiVL4y3d4rxO8q6IrIQ4No+
HY7hgIv8LiB+uGs7vgXsdFhWXW1gZZDK3qkdEoul0BXUxxgAq5t/9jqpxUPvES37
65IdD6O4hhbJ6YIdGFn6NMTlv9oMGmRHCxJyjH4cdxyGa3r9skqCCWEHpoaFONFR
DU0ZX7TFZi9nyjQ00lnQMjw4fcRHQtFFFnARcMdFuH+OK5x6dq6M+FDnEVKoS+vW
XAS3RUCSTZQE5DHHVYb2cR748BaD+cdbVvPR930WOfxJ4vXl/7KZceVjbu8seqg9
iHndY1TjxaLVmhdzUdQTPkAeyHFFjLdChYXVJjqiOOyk1dtB8CaNTgMEKvpKoz9j
2ZOUjaTCPXTveERqlf/4nou/0GQrq1eUjbMZ9BPHgN8xnHh9KOiWbexi3pa+eGqH
CIF3CtsKvhKTQQDya/Qr+MozKIBq0QrjxxFl3zsb85Vu/vIPzddyK7OVsvWXKkkx
ATLW8eukGy1YamFfS7ciiFO1Qp2TtmTm5u8bKxkBaAsLww9qJvGShpnXohUv3yzv
E90Ljz/mAIgmPgL2KKYIR5IpYXPwilNY7AKvV5LtujBg2qUP7qjFsi3yZ/44Irzj
Mk3mxNhCO53VeXM81QO9OB0A9FMoGF2UwJ0W7Y/FX2sHTeAdy2Hzo+/okOkNBFbP
NFPMm3wQ2/YFReDRKdzEs0pA/x0aDp4bpbDHmPXgYYKcPNLtGFMGn6tXGhJ4wl4G
7Zt1JpSONH3ineCt29P9+HOAVkZ3ALKqqyNBS9ekFESxXjKLwQnHZsd3U5a9txEL
apnQPmXRQw/1eJ03tz1s24dEN/zPeL1hg+jp3lhL/HcreqzJx4MqyMehCYYhRevm
tjmAeEN0E2gThXAaYq79l5zRLhqoH90I9kEb/T5utV6FvCMH0bNfMs1afFmol5OP
F6HB9xBEsvujryw+aziLM+EUZpFXW+hytAQz9+pxb3p7va0KUbQMggJz+diw3IxC
6HelM6CuBnD+f1UChzErKERjIRaW7vc1Uo9vGbsqPJt+bCB9a54zhFQJLTwcSNzn
KIYW/5SY85wl7tb1SLygF9D2UsAO+YxHGcqv2tqwqkc88E06JQ7YN8/ba+ib1RM5
c0d5Jl9HCvY3vG/t1pCbv7YDm5tM1+d9zv9pdkJ2V599aDG1SqILarCmt1+xt0bH
8owkLg8Q0//aYvS/i35EGhUqEAkvQwOYwK0XRz1EfwqoHx0CcJ//i3sCsJ1qCMy9
Y36i5P97h5gCKweQ8hTPhOSjfbQexTOO2ibN3C+kJ0VoXwPP8gRWWAOcuZbxbi7t
cWPCgpzJpAOeoY4qn6ZzOEemd0wFEJFtvyU6UF+u4Uwk4FDwrldFKCvOayq0Fm8m
ZzVLegjmdsfoZPHbHxPFQl4BaAJpcsDUPZmvVUaXb0l8vtA7T1O/kRdwCoGcxRWK
KlsjRXRrejr+WMSYrm1aURW8JXH4Eni3/FBYK020a+WhJUGUvlybG7X5z3CgoPEi
oso31GFVQaL3JX3ZcqcFVIUOMcmsRlkSIeR06qxghO6y+5QbFok+5x63cXDbrJ8u
XCveUl3Xr1qfAqwk5ZB1QuXV8XVlhCZfbF95ng/5ueHozqKQT5CCmxR6GO4+XyGn
mIAU2rcAcZiFIhvd1fGes3gzKCESgBcCyLRXpFBUdIdLomyu3aQHXQaIWP1BDQ+Y
xItQ5HEM4IBQ/kPdyuRKuvChkngKkcXYNHeHsQsQgkdtv8K/ptSCGCAj9CK+nKDT
8BrFKqLP3qRnij3cODQY081cjGVtFiExCLMJlielwj3VHwSCHgTJG7lF87egyoxC
rH+ghXtOIhpEnNsa5T/PJVNu0ELE/29ZnOIg13FWvUuUnX1QXb5Rh+0pE0oRQ4rg
5ghhnMqdHWgvHaExqlv6zMd+T7aZffWZvT06qmS2t1W1Ko2x1hvuRw90n90Lvfh6
r/Tuo5wODzrscfbqJ8tHMM8afUNQSVQAbalFpvPalBaL401EGyD5yme61Q8ZDXB6
nLqI24/VcJg36tlqXW3hoBefnY4yWm0LLK6aEP7DHVGbvbHob+ZUIWCFxsVGwT2I
BRc5B0ircmQgxbuK7i+yGyktA5a0pfMI+71C3DWfv7kjCp0B52IPCW5go3w8BMCX
48PATtAzQq/APtpS7tmEM/xRp4V2pDG/6ZhCeFVrbf1QnW0At+or2kKwppnHHHfA
5UwCTSmDTtGeykPr8s57zX5o7NhQs5SgDX4v47Yr4Y3rGBVqzdpU7QhhGWmxw356
dUwGVKwnYAf5+u2I6+OLaThwQrQk3MGaRsrhPB1WOZ7NvXzE/tN6X77WNbUPUDKc
YDUKQrbMAp78Y+UsM3bc2t87CmdEUiIF5pGXAjI/RVdi9hm+c6v2EyQ9NwMDq/1d
clE2GidnhJwkn0Yir+uxXBi7l/C+EK1yXX6BZ4hRopmjP7+iE2WVJ8mInPOLBU/A
TznGsxOw+hqODDnUqymtU2UhzEN/nGKnbgu3/ABxf6pd2ZtOclc28wGBjKRgSnHk
BovK4jpp+qU1xub7boNCdkiSUNG4FeEQrzaSeptKkmXHXgb+GyTAESO0RCri5Ndh
T7iEGQJBbMaMKgI9IPrx+Y5HdlKqMJX68eGvRoMZvppkpz2NXUIcbaWEwplODZVE
1yadsXoyUzuM5ksVcsv2GsdiZ9L0AbTQLMqlArKqPviaozyJ3ojgq4AGGRSICUuI
uBwsCxGgrMzesa+H75rzGM92J7Q770MtlaInoG4NKgUhPcge7kBdnFCqaZuKMpwU
GvcSi+w37m6EC45K3PFBHBQUetmTmsQCQAlFRxU8dB+mQsnMq3BQ7PJkdN1xKMcx
WC/ABOIHWroo5oJpwuSRZETQtvHi7KSbhNmOvGtvOIFAr8Z+R1U33WanedAsnW5U
CauCIiZLy91xO9xdaVJ/3BK+J/7ZGZYCjGLfk0DmsmEMSJoN/KRdTPKrzAsFhUY0
tLzX7cpUTKpJd53HLpXBPs2rUfmc4v3hY1TTU3HSl1aFwM2A2dyV/iUJOQBOCeky
Ok44hxTyWaRxM6qupINbMSeOVg/bf7vPlQbANGRCtHmRl5YyEMwMLv+C92FrTxht
NAw/kp+HYO+aFpyEKVyWylQQBDDZPY2pF4XrxAa1AbdhZ7m8SsiK4Db9xW1YMCgG
CozydlF+QzL8pUt0HPdm0L1+0MRFqxh9q4MxMPg1JyfVDChjFtWC+mKg3jn/jy5H
xznicYXIVR7ZzfJVEbh9/wJA4AIJhLe5q82sf5xqdzNY1Ns7/rrSKUEUByf3wR1D
2z88e6bsatXvuKD8hwRwHnxc6/wan0Ee6NfOh4oBw2M7BKlnGljsV8fVVazU9mFp
DWTphDtvHHQed3y0Y8IWg1ZkEuwKsjHWCKfqWGu2uSXR2V0tX70LLsWUvsiwyv8R
4KrGb2Io8ud+X1POWBAyGppGMyokbsDMLsUaLLtCNPk+zuIsi3XiDWm47Z66H3eE
xXyDX6xb0z6mi4VV5CihHzeFj0NR/8b45B8g98qlyUPUPO9lI18lsBQWU5JS0/1W
D87+tp3N9lhm1dVcMSQOJPZoKdgAfmry78P/CoK76krwfqkaCeu9fUedJVuEF3+H
kiYsyJ2eq9k2KEYUjg6lPsLe8MPYGbQziJ6ceweMHopQmKeDoK0GcossgUE+bj8e
sEaUmNYX2KWagDia8bJpnFniShroIKY3xXBiULULHAxiFyb7K2qw/NMLYwUf7NmJ
uWXIYj9ToUW9ZVr2PGOg9DfDcj6Fr2BDC1cO6zWSbhJWVbDS4Jhz19fODpY0sbkl
g0DMXs+ylSNZd7A5TbiwrCbwIGl364S4yG7/nz9vSRwHmdX4I2rELyZEysUC/I4M
HGolX+p18GeEphouWLfGeQMKIhBNOnOlQHK9K1XmPkJVUvFiSs3orrvW01oBA04k
Yl9FXxKQgt8K5Ch9iRJypkNsVbKWcjSMVNxV+ck4vFGeSNIv5wpE5DF/jNFnbl8O
zZzj7U+5q1QliW+onhOHKICiIVVLsa3ZJ7z0XicsqE0X9drTK4smuGYjsjQBOVAX
HAXfLd1vDWv38aYSn266BlaMZuw7RqjFDb+TVIThYQSU5eNfs5Dg4grfpHwnVe23
GALYer69IqqT2upx7RrzBhDFGhoUzUucMIKN50+Qfl0/p36gPdNKciITc/GBU+iH
fd6EqWryAc60lvFoIc3smPK/i2OuoSq4R3R11y43m4X/FzoWg5/5TCNV6uiGaLId
L8CMes78HQANEFfy7lCYcXlozcD0jbkWC9pK6elHx96aoOszRRZhnQbBMQDDhaeX
l1nm3hCb8sneP9GzOYzShdkLmvUnbVx0kk354bPkXq0OfYu6I5xlfyByi1oCnanN
SMfycHrxBS2nxvguu4MKsqz4n9XEblyRjIzxMEU3qX0SzsS6HnMVJ4dRAZUicR7B
ZuZDROyU26TjzjqmAvrkb2XMa84NyeM5EtEGBXJ9mttdchJfl4UEm6Y2W62PhiRb
s5D/3xcXvTEOiaJIEFv2eXysHCoSdmxXHAV+A2UDFZtaneA9QDQME0zwFpix03H1
++jo0S4iBVAAks0Xvk3uhF/OMClWFpn/NqJb2SIkBmnqJ+ZyHgtt0+rG8OhXIMEs
h27RIMIGVIolg46kpD/yGfRC1BQ/PxV1IMxtL0p8M9c8m8pQjegcf5JZBBbh1zLa
BZU5OdylmTrAx2Ae8u/a3edit5qBROh7bY+UfeYY78Oud+2anL9FkPah+FVBCVpY
EZwIuchl2AY0Uswss5VxEqgQhyUAj11lm627JlyFSm2Zxbd//5UZkAWLFfZnNRv6
Xb70yRcH7ImS0BcfcB4wN/D8xbwkhZMxMC6UsAynAzDSQnxcq8MPCLaxaemgOMYB
MAqrltuWqQ4opbv+vnFuUPWU+Gle+COtFnkXfGpxsoSv5hZkN9+s+VkCJla4I1IK
rN3fsJgF0UOYfonTil/I7JB2blWCQEr3uB5wcbXipQQkRPWWJFweLgfsUkicNeGq
J4vNf734hQ8TGQr+pn38szBI75VwzZxafb4DpBtr+hb/UAmUtW/YpIuXQzqcWhoI
krvhVmPehglCE5RhQCSO2MClFQVAu37S8Fjt/XeSPqQ7bQG7my64v71zP6v8bB/o
AuIRZdUGbEoA3ManXnxSP2v4YBYzxzJkHpsBn1XFSO/3qwgHM18VcxEmdxwDPO/S
YUTTa3w3L1dowRVQMXN2bjW3E9Zu0vfwWKdKQK+HcnY9+zPTxqnst6T7yQTqdlq4
HYJenBCqJaMJfKLS27+Kj4Frd2qg+NUiLnM15pHI7o03m4mG8OlDwMwitSfz01df
BFf/+FWW58jIb0BFYQeT1mZ2O5x8AaLpueHWr27De19Q3Vi1abaWWrjGMC5kaCaI
86cni/yiApN4VhXGGl7c+vDFK0KBH5so6zeR5eyQ3A6dN1TkWbInbIGKQVoQGd8k
x8KkT6wGzp6Fgz/1IUbEb9YnjbiB/yMfzhMAdNgesh27yZf7KzWYqsxHRJOWFrSp
SDmqpYRn4wu6N+7+Lo59+FB4mgJ3KEmuTzMF6S1KT8o5p8CENz8OkQEgAxkDG6Ex
3+98hNj+v7d/hN77MYLKvRbReJEFyUupE7NKnMl1wANJNPZ/P5aR4qlF6wvSkl1n
CzMqEz3tKVolQBvRshsNuVOYUuJgqfN+XIm+AwlhJoLNz/LfQIf/ai4mf/sE5ySw
LSRgqQAuM8WvRROBwywYDH5GlI//9vAO+NsfOkVpvKQxpON+my0p043YxpspuUpI
ZE7rmD3/GBgPCWnRC269y9a+EL63tCv6qM5Sq9Cv0FsosA+aDimfVKfguz3eIm93
/WcR0mkspKR21QxMU7RMuHxU86S9z3mtOLj3Fo34eh8JbfniAqpdBMVTy3cJGoZX
h203hfZsZMzcfy2ldKiJ0yozu4aURdMOMtG0+UekL19opXDrvTrJwqTzArDJ7oxD
36JDR+KkhrlknLs+7/talNpvA4mGjhqV1nYSnp+yQEo0FXKYKB3xMWvK6sJbbCUp
at9FW4Hkx1nSTkwsatW0NyeHHJtcZSImWKflNsB3UUGMTiXx2j53ie/ApW3FtvXG
RzAz/APlWyrohdxGysPjg7Xr2gdnpCVckh2KE1tQKpJrL/le4gu2CDpFi/8XRmUb
eyrLX1DvS7fXUybxXqwS2UhI9+0BrAkJxqfnadI39u6KeMf55SNq9GXlZpC8FUEX
lhVbiicookuMqxjbIbivTCqz7Pf+ltQb60Lbb/8wzf6cXWzIda7g0Lv06D0beEhL
Z4IpUCJxFB7UPd81eyBm8jf6UY+EGhbzBg+eVQa4Ax34+TosWHcSRWzgkJFNe9V+
Wz8cpO/yjsghLvmQsOw0zSN7B9fHC5/IsmQc92eAHtkVcS+xqG6Shqv3gCYAFNvH
fqzYErwa+Uyi8dYPkiBXiFT9a8jn4b1Xu8y3FBNx02rvKqnRO38fxA6FHPtiS970
cNvqjcuKC/8bEk7owbPn0lVUdgRXlnIFltQYj8BhY7D9gbIObZpo/+GQ1yzxWvZc
q7W9iWGRWJU7if2Upo3SssbBTpS2z6b6qkmofJJCflWnAonN2irJPS1jE76/WhqK
tuBfXcOgmDa2r+8Xoi3QsHNmoeNdCH6vUcwCWgS0o+Ny7vWR1cwzvGJnXuzESo2N
/CvUSk3YOZwNp9a7/WnLRt3KaRoQGZ6nkFnxOqqAr8JCjA7t9duuwpn9ei8YA1aA
kyeTB8Ct9OjQbTrz1vvf2zUS0cWNAzJRmAg2AJxcLH75db4gkkey+Fp3XglR0fD7
EuwMQ+xO7Ho0zwIuBFEKN3quhcxi2RI8M9Rs4OwmFxNexbTGpMdygw3aH61IFJXI
C9IV86p/Zyb78LXAjC1XUflnA/amqasbUDyOvFF/bSw/ylT6hroKfnCbd3KiLEtR
pPlh+XR/XJ+eeOVh4UjR9eEJ5ijJIoXzqkg8m2TyKXFRCjr0ZPsNPb+pB6YJkFE8
VCMFchwOoJS8ZAjwn8NNX9Xt0OO2fyatkE9QF86UZWnZqI/jrAogLlVZcoZ3pP91
2lk+jDXO/p1EwN1SAx13mUuCqRxU7OyqDRtl0bPSUffUwkmux0Qf8w95WaivRnKP
uYGuu/Slkl6wIk5kyv5LVYFmyg1GqlzIfmbuQ9dO9H3O4X0A7InItBj9/NBH4xT1
kqGgBRiFnQka/EKXzDvNWgzjKXZXUXRI7dMYzrmeV4ipNJ6RdgxYqzZPwUNnY83X
oum5egKRr0rdaDXsSV5tns+qaKzoOVVqPJNweDGjgJA/mhRk8rcXedj5IuiZSYF1
KnmAbzL09L2gG8xs9U5I47cNC37vWc34WYTT86PCH3hjsxZ8qESDrU+bfis8roXJ
ksyLRXQTQGOqQWtLRG+6UaCJMy8IUX89EVHld8SLJs4Jzbi1qTLB16/IVA3yN2jS
i2I2xSmhloXdhEMRtMfWqk9ffYzihL7oM1ZbUtBws02uDhLz57x17IZ6+wXbbGvV
fTwfP2oYM+SWCiUstz8eZpnsM+TIZUg/NI9F20M4F/OLBTB501igyuU4OmWnGTZt
JFoAWiytFYEcMa1bi5+qjsOWOUWaHdy9Fj4Jio8WxSCYu9U7nEC4WZ8YxWqxcsOo
eXVm6d7VO/pBq+MntaVL1ygRp01LD/RxsgE6ucYIUpLegVVWE4HbesqDJWktC+RO
lSPlY+X6WMt46EGDadhcu95M+Q1WOkEXiuEKLDRORRwrEvTpYekhXJQZ4y1ujiy7
BkDUBMIgs+76hBVDn0VlRt7Jh1rhIOht8TDnGc1mbWB17L+E8xmllpbMeU001aPt
aPo2UU8CAdGHQbPn1DQv5l3hyz6Hydm5xzKCCHr9CitGLkdmJYRWR8VqGjTi0dq2
Tnk2ycVKC7FlEUDnvgoeRjC5hstqo8Mm20c+QRwjMr7g8KcVP0RqksH8VjrkZlc5
acoSnxKSzgp0n+sAU3PpijBqMIFOLKRtB2bdvjO81xYdUmqAwRSi2XMeSOBH/qWt
aetbEsYU7XpNamXHA6AFkd7KUryK3LUZZtGwsgXWIemGl1Ppf6XIbIGsrawbrg1b
DLdZnKHDiZmXCXwhfqa/+nHpAX+rMLiMXFIe+huYKqJHaGyRi7odfTF4jLTBIioZ
YIX02woEnA6wlSsIu3jZohd+bxNkUxk98HFQUfPGHFrC4Rsv5+wWuzLJbp3A+Wyv
VPr2PQbYrUqz1k8xy6/lvfCwTP1SrWdVbUZII9Mg/b26V+oDfAsXUPBZSZ6WwkFr
nZg/zZX2IlSEzsM+27YKTEfvirTq/hvmAP0hoVx1LGI/SMJpbCuSYr0grEfLuan3
/sDWYFSSjQxujWP6nUgWdS9T78ryiOVVSyTEFtEq5FEhpGbQUaIetG3SlxhQfh/h
MT32x69ii+jNK+CTmCLc9AZ4DjiHgNB5iWW5NIDV5aVO9IDazPSwQNi6aKBKNkf6
bUHiSxkNsN6WvkXjjLhRWyHeQu2paiZ4CYJ76g5aMmGwQX3gKGbOwxPioXX8QK4N
+G8SdNOe086og9pTdRRR81xM6a1UGd4QCR4KvKog+ERzmjSWu9aAeUoZXEK+hsoR
lsHtkWIrEIan9dwqWxZ+Qhxdg1AzfMnf4TwZjAhrUnpisJ2ocSS0vXFkEd984Mit
QjMUlZfyWs+Cd+5GxdrhXEjmItIuPYiU4MKy568sFv9AIJuZtBfM8Ry116YV2QTV
GDCayDgsEHUQXq5bHTKdIBoMC1oLKspaqRpsyF0kWVFhPFMvXGYjOFNVohcC7UAo
UhtbsL+JkedayriA4+90yD2kPwrc9C/Si97Wvx+d/BMgZgYORgeKJidVpsiqf6Qi
z83zdyzeBruBuqDYz+hPHc+iSY4SXSO29L9mFMdwPqdqlujdMprFeYDwHWJGpPuI
djy0wDNTJtjHdvy/7wWYveq/dHneN5Td7cvlVE+t5OCJtCvxl8eW3NNvT83QJpPz
8xTRpzOwqGvmmBOch8Zw6JQH3EZgVKLsZSd8l2b9OLcteEGQ+QGP03IZkOq1h1Ku
rrPMwXFs43oeEET/JGSC5TTHzXMNdkxSKP3jiap3Enj//EP/sUgfKOfg8aHjVn33
B8xjErUELvfNk7d1P2rOpQmjra7XaBDKzSREAkrPwbMxZOeMw7Z52wEERodOE9Tf
eHMOHqhBAv2pFXERcbpU/0a6OgRg7gdbKVQAG/F2sRslojyVBvFTZ+Q4gdFlSoZF
RgZc5LG5koL5caukmKzgMY3d8/xpSXB/d0Wrxvkc/pVkTNLQf6LVqOhUru1RVQDj
0e+6Ezbdx3TmXynvOobJxnhK7S1Vqg2iAtYqke5J7VKe/e0EIz0/llAtcoR1clwk
3kvrkpDFOQNUmsPbCk4XOoPgSXpK5eAy2NH5CywHyOfqC5Qf/wrNTXp1kcAWMyhd
ymmfo6SjE8hR9nq6njAb/AUaGLN0MnovkoXtVZAFWRQzxgFjE5lDxNOMHi1btste
QDcqZr3QiX82vCLIZh9y7A0qFD2SmLn4u45klXRmkALfLuf+B47a6ZHljtmCPQ22
VtvyHsMV/iVvuq9QTBcgS+qAuURLzsI+yKlQ+Zjj5mtfHKN7OaByJW/AJSPL1EBz
EL89V35/kES1sxLrK99ZIHIfEalqqNDqGtzU/u6353AqSQaX0GST1q9diC9fyCqe
7ikpwgcYBDO6i1gkabHoYujiBHmPkkcHFtK8fyFkAaO7MIEzvxfOVrzHooFpySpG
DXwvEYig46MMBTTAyzmEqJVyWcgBGFPirYPCPDes8sVbPq2tJrCYpxRQZkYOC92e
jSUvUol9WSpYL4u4Fm+7Oe7CYWkfslglljyTVASnhxkIDWAynGB+uDXDtJVl8M1u
aKqPXZ7tBbMucUC1iFXziLfCz9/SXN9qZD9sJWNkw407qBpAg6XB7B1yYlfqIXwn
1C0G4d4I86BKVfAPA2BiXXMXEZDnSkZ7wsfeJSQts5W1n8Tyu6RBRLBCBmYZuxvg
9Lg/+Q/WYzTcxrwZDSiqvn5keCda9ERimD50jHagEPaj8DQzP8Rlrd8PVJW5klep
YKwIRqWhy1T636shRTRxAT91CDy2sAl3loU78Q2YxNu2mqAuIqkClUgmsE5TEl5r
cl/OGBCpvKPO/RbDYkwpIutvgT/bI3ADNdhYNldVQ3oVhQy1JaB7SVnuM2rfR/0J
F6/GWHRDFA3D9R30sa+9gto4IoBblVZ8dsJU1NAqAEWmsWX2hk50oAHbbnYH09kS
66Ch3vOCGJREzacctmAlgQyqPzpDmGzEC7Lyw6Mo0Z1jxZTVpChVoOEAJocNhbqY
lt80VHju3aeOEbDJGTqK9Yr7pPGo2eGgK7zQSQpSwzdi3Ef1DrrkZRitR9pzdrAT
5gmfZ9uGmAZ4IVqmPhELdTH4PXtrhL4+2loXuVjZ8PtDnG45g9kFHAlVGg3KzFhz
xbe3ueMsvbc1VVDskFmK5uSmvy25BxXai7C0tmZB+J53vk+vRPiQAtr+7YzxnZV4
/wPsW2RVbmOl4zkd/Hyp6Frl00+i/TdTD/LiEJZpbX6etUgOwl5Rlb7fkuaJe/Ds
Roz/6CGaLpLceZgOnk72vrOJtfmJU57MWFSTaRCD5W5CQdMsT93+x3ksIUgofdRH
bH/QT4gLHm71ruBe0sKuaO86V84szMAsJ4i7Q7ajWinFWLE2BkyyVQ8UaUEof6Bb
Zlx/nqAlGvEjBrrnv1tKxQC71cgDaztXI7hkuXaf1X6PqHwtSOSXmKLxAacM42mW
WYpnmKl5lS589k3RXcpu7BMs8nWWlzoA4r4oJPlN41Kz7YhS4AqED7sh5gVIRnNQ
bgFbOfwXdS5YhSLCcBOWiQKnOpHUtleBuFCwzxIiEaXttgjLup+Sl6uS4M3nfJii
z92p15cPERwZQ8dECNMFdsnQpfX0PfPVNhnA5gbk2i8YXmqsrKwTi5XBaFUKk+yo
rrcM+smopOC2WX0NkbmaWTymoFNrVQl1EcuY6Qdq1NiOLMuRzrnpnTuO7cpKkHn8
vhLwnCZcEV1QJv4WejChJs5yKgtYp4uZTjj70xkjRu9n/Rflq5tv9lWn4f/GiyyH
UdsU3UIEMWdwkULTtHAzf3vYCkuRNXcK0a0KfScTV9QuIj9yzpo+t4d4nCvfq/ub
Ek/FMNsEcwfDraFsF0MS6GBWdNZGsz7a+FFGkqbi1L4NYWQaCq4OVvs9+v4ROSl/
WnNYUW93PGb35KQW12aUtCcfbbSNY2Y3KyAQSDUtsUjEM2hvdv6V4XbldYqf31qU
7y6MwQqU3H2jzPSmNgCAfEdgl1FwzCTiwxao1ipmc0FkoIp/PslyJuokyP7lY1T0
gw+Mr5qiqKQqWwDz0jag3OLSUz+QkjlHo/PwLDQ3wzmlNnxVH4eImBF6gKiytEXk
bB8/fCUDPfL1fdgL41UTWSF2l7Bo6SXpeZuSbawAd/+frYf29zUzpGvWMZVD7A7X
pHw1NnrzRyV71LNv7LPtOS896nMz+1ov0T3E/J6Hr1rVd+t+PJt1YEluZcIGUVc8
vH9wQ3sJGnadDom7eoNSh0i9YF6Vu6BER8wERAMKkn/KA18R0LfAyv+Bv+tAyjgH
ZzuoTArnwE+XvdEl1DQebJL9RQpXkjWuZFr4KT18vYvlGuLImpJsyxt/76dcIJtG
VBuy/crfKjHm8ZSRc4O+czWWCRDrkXbZL1hnM86oegWTJY9+8vBvCYcg8GBILbNe
2/oF5cqukDlcv+oA4MaOOaQ/dbsXzUiNaERJx0RJgpnzZz49UyO/ogQ6lKI4FWTv
nbcusNNu5xcnDRak64rCKlOGdYVC08CEmCkg12zQYLrpP20hY2c+d07hebqAe8sR
Q3IeIzbyUVXHAP9r9Or/CVCC9QAYcGjJnK9qOvUVAgHfeXHL8QeZvkCtJp6/q5/M
EELYxJIGQo2mz1hcszERkUiuxCQ2ChQfy4jb34HtfE3z1syRw2uSCmJsSKUIB0nH
8TvRUuuoecf7b4ziRbiyU+pYsETSPFwvW2kW7mS2laqgIdZbQzbAymRci3cfdwXm
vJbOT1R5QB5vLAtU/UYX7MMWf9EJZpkdaQoTBnqIaLMnIqpuh0r4DaFy/4bp3R/R
sEei3gKxCyWsW1/H8wi9Ja6LgPTl2u3bAhAwcaELRug=
`pragma protect end_protected

`endif // `ifndef _XVIP_AXI_LOCK_SCEN_SV_


