//----------------------------------------------------------------------
/**
 * @file vf_axi_sb_func.sv
 * @brief Defines VF AXI scoreboard access function class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_SB_FUNC_SV_
`define _VF_AXI_SB_FUNC_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
SeyKGv4jN2EIHRppmCi6+Qus5MqzFNwDgRaf8Fh8lBg0c7ioaIvE5DJChXBPRJ5d
1fRt6pHzT47qHpAeMslW4Cl+aCYbP0R7ruDVrClv1dIVSzgDIxpTPcSWk05MnUHp
QSRdLHnfHphDrbqDGxO1Kc9aaS4KY1frBISMYMwQvQXjhCk9f/S/yuTAcSqeMEBB
GxtPWd651Ka9BGdB18yj9yX2/3AKnRvkKko5NjQjrotNlDNXPymZe2bmc+NPaX99
F2q1BIdiVs06jTXsgSdp/2fYBQ5dewkfrP2YLyH96AjEOtn+6hYpQ4Qj+v0y1jmQ
molguX3UNjEEQPfR+dvOfg==
`pragma protect data_block
H4FjlrTqicl/ukkbS8mXnwYoDPCiEHQp5ztb/B4v9oB2KEpZkFTJ43MBBt2yQIRw
vHdBSfM9lCoiJwf1n7Oks8Y3B6MZjOBUEDt9lS1NJ1Scpm3FBn355xOpIeaAwnCx
skvAjDoFfkauRZOEL4pV0vlfaLnU9Vw1duXwTp3sIRXa5Mn3liGxCs8yta+pXxeF
1xXe5DM1WRdaTMgegOGaFzddMlRS6+f9hARH5fun+NfpaaXnwxETIMGa74V6wrtf
BfgYCiB07RHHN7X8deQDusLGcFDppfNPggfywj4l/DXQI2+f42gU3FNTpwFlhDJH
HHI1Its+9ugysU0x3czYpLnbwyIl54b29H76iSVyDR2nHP6lPNkVZ5hEB4eOERr5
zlOaKviivtawilmgQpt6cjHVL469B8/FV5jDTDST2nCcVgHPHOo7V8dw/gXYc6Kx
d7fbt/83r6Rn8KwstfrybH53uZYyP9cMat8vVk8tQAkYlLHhrTM6FQhtnz+GzVmT
+PYM8CVAcOdq94aDF2dOciXUgB7zNyWt8JVo5Gp0W0PYqPlxf24oKzZrQ+s7fxis
9M5ZrlrAf8A5nVkeX0iJ9skn6wsmkgMPRYWBkv7wlC6GWz0O7oqrJIDUvna7GFJW
cnGZR4uKPonV2UNQz0rcUURQxv/Z2Js+rrQ+T1zNB9IR7bY9DcX4Llo4MYrEXvw7
e+i4/Ah3KOyhhJgD/p/A1mMTajl542nCQVkGd4XSgP5kZRs2NVdnHu3iGDdJHFAV
dswYG1/NKjWzWHriYZjHdiAlbIGX0o7OReDdpdJH1YaKR8l0eVDAimoSTVnwWpT4
YGHKD6AhcrUKffaIYeRn7GPhwQsVC8404MsIUdmp1+mxIeoR+21A7HHoJYCrP5W7
Tdd+KFnYUV6mxdaLvaEzvthUoYwHrI6a8EDE8C1CgrOptm1BG23K90vkLR646GZx
YkytH5hyw5nNOYneNrsfKN5cFSm1nHKEh1klbNHH4cL3dH1JC/kdybFHdQrm1qmm
TBNKx06qyuNt8qNpTbF++151h0cTUi5WDIgONCPCAy4Y2IW/03Uvv9XAFookdYy/
uI3YGFcye9qDFpO/GXNCMRCig66TmQVf5Z6FaMam1gpE6muH6l9+c2OM3v2yefHh
QHeuq/njLQFfyaTBjgHkEv4f1ggV8272GxYEXlQpsSNN2nU5ER/HIauzZlaxWxez
G+jLCpSJRHaTqnTjA7NpnQpl29K18v9hWZOqOyl6/LZs04DNBBwnL4pSU6+b8dyg
phZHWLLFLKRC46b0yU/JEVCpTl5JqdybwUlyisU/rts8bHWEZTRQZnNh4rA4Yv5C
i0r9QrO5xi94ydW8HzcBP3WZmYzxhKqLACKu4RSXLGI8Xp9NKmkDMktgAK+zNdo9
p2oNLEQEXo3TXPLay/HmMKg/ygrZyJOiZ6IhLNrOFwg6CtyciAK3HRVe1hTNzrC9
0Dh1QWiVYyL9TVqyBv1hjziqF8JS+WJuB5L1fmLU1z/44H4e7fJ+bNbMXIbdHQIk
XWOjkbP6b96GCeiBuCbFSIK2sfDxhXdAFOMz0AiJRR/Kg6+7VJsNvnIBZycGXIRj
cOCKYrtQtcsKAekt/YWWOPcC04J2P5Z3RS0eyz3FscKTdicXm+oeqyhAZ5NUFGLb
rIPZaT9PWKN2PdYxPdAuC8Yl1XbvfAzuSKScZb0kW9nXKvc9J+WmCe6octdJhVtS
AM8nLv5x2LsiFCs1hqVNDaXR/3TKGgvgCx0H2qry0N8NUQpVOB8ej1wkk1YFNS9n
HkzkRyN3rmVxsd/46O5NZGa16VrM4jD1EksvJpVM2jEx5DKIeYlnHpZr2cssqTaQ
AWqZ2CCMRasa80rZTlZRvEAYa7DSqNnXXZ7uOKUithMZ0f4F7B4VRVA74Kg567Iw
4IPkZtivWmR2OqWQVLcVTEvJhzV6APKRWd/SKUaEl44j/qg1k6144L7k2JnDuih5
7gOkA5yYZyytxt8YG2zKcZ0x+Ed9Riqc9cWdaoEpRHcdVnzPeVr5194eu8677s/i
AQvZWf/OdUtkZDsvAI5Ml0OMaXDYhAsWfeLXh5CnrWuIRhSO7OrV7LOf5i2+mQGz
4bwsnkRC2e/dEzr2Q1/RyHckrDY80RS/L53wJqcc7AuL8Xn1zEWp2YIPBCsb35pN
/oAtaapdixItPqyGdzOkOSoi1l86rvtUKTLPnt1Hm1mMknGKZtjeRnGh/OnlbvtI
gb+VcJroH3p6a3qEpdBzOAG0pr5Gxk/cLWFO9i9kQqsVnSd4Qu5frVt2dJde/iIT
SOXpUSTjhdy4SQnqrfpfSky3RXF7lxkPtoaHyn3PqN0Mt5wRirlUAg54yz9iuA9h
QC8lTIizQ0WPrWlwk9RL6aC6suxdu3FZAX8bNxB77LoetLnZiDycVXGvdpU+RAzB
/DWNgt2tjbqOznpTvnGjtCIaNsyxIYwih9YQM2C/rgVztnBt1S7tBj6BHDVrG4w/
mCZB+sf0Z0GNHj3HZ2tC2EGD6LcEbKYlt5dzjyroBNdYmuGSsO37/0NLrfSbXq6S
FsP4VXZxRJqQ1/psRm1Qn4U92p1SUbVrRRlJtkROreQMr0dUjQLyPRMYutSENovZ
AvWYHZDmd9YY42a341c6c05ApQULGYHZrecGXtKzUA7piczJonNjjlu3xs0BGvYJ
4VbzBSi2wKPDFakh0QYQfo4R0T9fgAwhcyASwH/Z7Wq26qItPfoVDB1RuV2oZLov
0OiM/gBGUCGm8Cc/3e8qx2+DST42rKGw9x0hs2i1YWYgZtF6DVqaBImqCwAcghYl
4bU2n+0Pexa0Ai89KC24j8Zwiv+/E46rHPvA/+/Rhjh/WqhKFfeY3eoNTJcl3lYi
HI0zRC/Os7Kn8F6YQpnyzhRUe5hmd15a0Tk+pgG+lpSJ/wPPkDkC12SlRxy0g4X1
xS6dwHXr8Usmi7LTHOs9p8NZL3lkwJaszdhgyH9MggL0kQEJjEWsL9N8PdLrymbL
b8Obin8ZhGZat5gvzmu2KSc+g98PFAMcu7T8Ik4XrC4AAtcVtrMgbI/QPZoeY6QC
VyxxXYOQz+xAWzRsGhsXfQR2AxPFQba5X5Vl6d5CBjh9T8wBzGTe6H2NyGqfn+PJ
o6Nk+SFpbgCUD3ptWc3OIBvUFIe8KaLGhjknVbL2Cqwm32/J+Dhx0NvZfkV1BRfn
zHVyxDlDqiHrvTbJN4Nwy4HFN0wl4+T7Ad0zIiVa5vsGwUn5hKQEmXxFA4q9GlSY
aIVcmY4Ae6U/EB+cmW1H+OTDYom/tKLPKIpLdVPfOpAgZUMekDISswXPy/f2MFM4
AJfa6YEza11BGPeidyQAGtUhGKauc9RQRptv71AZzEAq5hbreg5B0RU9gViRclv3
5jtz2Y8XWArfqtYO0oojsRHThZu2vMIcdGlWOH/PkUj1+py3DBO0+9/LXhbys/Hb
cfdSjhgvuNrtYeiarDY46nxuedHEhXp2bf3/+6IFQrfxfFd+I4QyWfKDOVvuBMeS
9q9nFtR8Ft+VYW4qVL42ScuJVnXUZOOhfadiUwHRsLaZ+oKlLjbv/FSbIUvXm6UL
S1xfARK+9STIM2AlPiVA8mYwiHLEbOEp3g7D8GxD/Axrl/cVdwYyhXCOjjWCglc5
g2FYZX7v1yAvHcwtgvdYF5Y/BiJhxMs5iWpIe1Kqgn+3Gut0St449IgE3OqzCmUz
M+hH1TRCMCLtaF6fnHOJ+XT3DsaJiMg5X7+UeBEUpNDpGlRXdW+Hj+z9Tb3yVN7T
tQbjdoOD8Kp3VCOZiuQyGH0RcGRRZX0Px+4+MiS1JbcD1El8Q7lAaHN9641QAD/p
M22kGMvICNyOmZJcyoGtJi0qQ7kTB4TK4CjQL2mDmn9YeQS04Um+qqux9rfKx1Pm
oXPjynLCT9Fdd9XvQPit4qxhJKH/YBS0vRJ2oMhJvubQB71uiln2FfQGPBQFaGPl
eKLdY8mzqmRf/kfYK/d9asBUrMxDcirSYgtm2YA32J27oQYIOXdqOIFBulL2IxOC
hWQ3S1Chj4paRQUdulgpEvl8/hAQ7VlMN6Up2btKygFk7aSAGmyfQQgEL0EFo86n
ZTL/f9XVTI1iFAjR2LruhSi/PI+qEGN3DoX2DjqVxNWIAgS+liekPpmSMfHcHh8h
u1eh5aYUOt0KDMcf8yXjIK+n/V1ynUZalN+YJHJGLMFWVAr31kC/bn9LSP0MaDZ+
6Qse67IxCF4DOJ6bi5EG4HuQEsksIP9iBSZAAulVeQ8UccywLxg31NN4w5J4wKxO
LbTPP4M+Cgt3iapXl8b8nzhqCImMRizaQM3qA+cqI18ncZY+rrRbgDXOJ5NNgWb1
0Xrmc7jiKfz+ZfY9Pjq+3iFMPJ4IMVDRr8nEwkPYsjWBrsJeAVI65okmviH4AMfZ
bTOnLgBQ3txixq7j42qdkggUXLw0GRYKqUBxlWDshPI4qBYCOOJvagMH7m2UYOY8
Ivrw2QuhssMpEXwJGx2/4+zdHLOc96kb3XkpOQHKWkgqcjpH8//adbXEscvpIZ1s
LEyLegW8cww7Fezb9b3/VWQESnxOsy7lY9TG0bXljNN2BVkjSf72uOBDwGhhnCEK
To6H2tHGMOFvFf2jOSgDNX42iAimQDvfToSTgqJ2trOhm7Cig8gWUEIeTtw+LuwU
jh7mLpgpiYpzfnu1OOvnSs90ZuBlJk1Tu4UfrRVNlG14Z3igsbFnfYUmaVoLkGMM
HajwWHPWfHyN1HAmyLw4mguMiPa0b2MSF+O4bxp7nILZen5w+DzbPA7WNjyBEXTd
+6DiTx0r/bz08FltWWRBNzAr0oOqxw4hsNvJt//Gz1ox9TA8KgshBt9B2Cf8fsRe
GgY/yJrecWmwxzOnPmiwpTKQCb+g4RdDrSixjknSvbElZL6PTJ3zJTx4hDqQNdiv
GluGEqDWx+X+HYgPBIwmE62lj2VJY017n3Unp75tcUtt0YksPQPz18NKoYJXfTu4
7ACk58UfsZFzy+c6HmSbgXIOWPvmbQY7YhB/QLCMO+eg0XtKJODKU2nWVSxyabQz
z8EA7J35lYOnLs9Oqr69NqTaImwB7RHkTiTJs8ha8vy/l9Y0/ey0DD7c3VNWskFc
M5d7MmnkzoCBbMU7goY6+b/Z8B8Jb44m+E/3Us/dTjFclOKxQk+CNJXgtUs+sCbB
i/WBq+ExrW4X7bIvkpMC4JulCUW0KHUsm+WJn+T0kVvYKDjdUUCv9rJT6B///Sz+
yRbcK4IAxNLJwsYf3/ULQl6JAGAqEn6ixfAvkFc7JcVo5plK+4F02f3SmA14OhSy
vNmYKtA4z0YLCbmGNbHiwgVx5RyOkPac9QbyaRQ8+AF4M0L7E7VPIPnIhMYajQxk
gK0B+S8scR9h+lC6uc5EkjeUujDJYL1Mbg0yGqmwB1FeRdPXab2Vkehq1lnCfCLQ
qGEsvznL3C3wdgE7minvkhtEcKiQ5eRDxHycu6SIG+DPp8Cj5Ui1uVUZMOho3aAw
LXQTCim7PMZ9cJu2855OFV1ntkV669nGZXeVZrHv/f/vMentYRtOwsEWX3PRwoO7
t3Hh5fJdKa/CJcI9vpFdA82IUHTJVwTEHmvkUxvPXzO2mlcnjtGxo52QZ+Av2CX+
Dic2/gja4JzAxuQB1lzw543V8dOI0B0iF3Phi3NeW8VmY+TjZTKQSvEUGTt6gGHc
O9B+FblCRn93SE5v98WsIGCwnIYHwOOvAcC2jH4kl1acdUBfmYjimkpAXXbkfv7a
lKCrpYRARlSM20JETo4Ncoteku7hC168RC04wdiGw/4ouzprVAdldVq85qp+3yP2
tPYLz+GO40IgIFO1s5PQgY0fHxeQfd4ZLGkDuPAcpqhuktCV6HXjNgbn8YHosBv6
0rz4O1aHbXUUHG7hAgfwCyIRci+kUizLdrTaULboDIj/aAYZhgPVydpJQFvA+gVC
oWz3hqqI9gwkcDP4yB8qhEFOccBg+YfLmZNWIzf2U54LaaO4KUiuKdX9Tk2ABbuD
zisYrf6xNbtuz5LWp01MTqwu5FKcFsQXM4obQoEjS39aq1HR/7OxvAiDZBwpSFZC
lcmRABgOCa9lUvbHoyaJMkx8mUHvA2/yIEbXbwlmoK7ivdByNRHe3jSlD8OV4Y+X
S9oRLbIVQHo2qR48R6kaCFrK3SuPxf+uSz39x5aViuGSpEbDE14Wx8eJqN6bYMSI
Eb5tpedgVJzaR2d8lGIaRUDoA/oiQihzPUudOhoAE2RLJr+LxOVcngChzmavH6Kk
GNOS+iS9oosqviPJ9Xa/8txVYOD8MqCAybSZ9BKDYUjkm0Hr2krBXrmY15iEr7cf
opjnbE7H4n6PirJ2QoNgnpRQAsZWzz/B99kJQkMY2AiZR5em+NMXW/MOtBQSrP26
fXwXXRb+5mumOBOCOGwgZ2HmMSWL/vfrqA0swZEtyzX+HSCqEJIrDOq3T4FJZ8v6
fvQLRmH6N9k1ZdwC7c/u7DqGI46JUsOZHr6zdDP4qmfB1AZ97tDWIduwXjGRe/TU
wXKFgcCQR4rxaJ9JcZfLzrSQHMRwI7r7ShFR6pGUfNK+wo8hVDekOMLGsqsgvjHM
bdtqf6Zl4hWK1V/oGFWI0amDvHZCXoVaxzidiIhoMN8tSmRjwj9eYpunM4Y/1baZ
RyY1GkiJm6U8JEKIy48p0YB93cgFEuCpLeFbuxNFt+QYwiLHCUhPvlMDXI0Atxhy
6KNTfuaWJa5KVstL6G+/SMj79Ak8LR1U5r5SMhF/RKmaPm3j/LNnZTimAEFH8AP2
jwLFdcKKU7Cur3XjyfWptqv0w4xcej6SuKNssdgYpTy/ymi1r2eqbqGKJEKpIEaz
Rlj6qhL1/kKiVUHjy/2hJGkhEcG4oi+4Ew5uFOzU02ulY/kzSCmmaAYm6nSFzVBg
SXXomewUi5zJBWtayGoAD0aVPqNoSPrQ786IBPcPLGipqfRe1tm8RYNCfCtSDeSw
iVC2+kjlpNleDWvakwe4E280NRbrzQVuOduQzo0TSqoP+r92BprK55He6yGTJ3FC
d3/xHPHSbuTWdtTyztrLdNxWF+trzooFdPTLS9kVxMD99jEfWNummHNe/w6wkCVT
lphyQ9LDVd/00dPGbbqfU9uMQrBQjX2D2tEcHnjbPUPrubb/XEkirwc2iBncEvc9
s5xVLlGYYIFQy0UnqUU7U8OlpmB1WzkmA+UHCXwznQXo1DamnkRuh18fV6oNl+Tx
+rGV/dUVy51zW4Mg3xCf210PBlG5MxY8H8QyRiM+btM6Thrr3hXFbIlnXImPQXbR
zNcWHWNt0V+e81AETI9Sdb7zXTQOMnr+yHXUIDaxkN69zdLVPVLO/Lk4aDZu4AjY
M9TAazwUZbWzkfSfzhRaS4l6iXd3wFYl/HfqQFNT5tAL0dNDatWhbl0sZkRSPSAP
Ba22Ww7/PD7CGV7+NNVX4updTLNtLFKdvM0vkTCuyCWr5+gtrO2zsqoB3jBnOzPm
gbRAWUCLACw3Fc7fcBTlsdiXOQLRKrFV4XD0SWMTOBaDeDT0/24p6941aL2qNEhG
TaKt2/ILPuGwMl4C7j6WYE+EmlxhfoBx3IRpccLeQ0qcqTid0Qi94xTVG4dxzte9
VDwZFNSLSxBWVgyHRzwURU4cF46zw+GiIWG1QqkLEe8ku7KSQldPQ7+qbTofgqAR
ZAOKSZft6SlSGI20b6HdMqVZ+vvzbp4B9AJlg/drfp9hDAh25ydBncnCeXylhM6e
eH56jsmQtFUfBMxyEbhDxV4GN4jw2uJNycjbGMek1tvCB2C7XZ4KJQ7T1h1FMkrX
D9ysaAqqSfi5O0rc8N/W+l5G1+L5ofyEkQaRMoT7fi2BuHpLmhnXWAPGYZqM61lj
7rfjy8S+ygHrbGbCCK0yvQtyaSIiwFnVGhAMXVPWeImIMDK5INFdUPQK68IkZsU2
SYZV0EeBgoFnSFYr3kZsUjMI3RaXmZRSJ0EOlV6WctmvyUuq+MrxWsA5iZVWg2AV
3ymrDtljWagIuXSvArBhShjhipCk0/297OyF5eXAwletuljuVgwHmAUxqkj2OA48
Ow5wiuX6b39/zDWvwA3HhLpvwVJz5kZC8dqpfvMvOMkg8mkvIZ/pWt/sbAm8CAYH
cpPAS6FagypXpNwnVgfjqS8f3Bp/kWFT/W/LPOuDoXzOMOgaf14mUswFw7BUV0NN
3TXKFSEEMsF5WeMrJnvsYC8BGwEUOSKX3CDwuxNt6NrfZ+cyFWTAJOTigyA9W2Nx
XvxrGVs0Aat5bKrx+XU+g1QLJ5bV32sWjbJ8bI5isp/hcy0DHD+XGYEBTZx3hshU
TDyIushs324fcCziB6YUxL3D+2g75q7/3Yo4QUJ/w70ByRCmowk5LJQdC3mr/DKU
+35LPTgvOUNyCjmlIoVV7m0uKAlC59ek3TTpsD7kSk3fQgWFvYDluhd1g1hOA4d4
nO0XZ6fiWk+6FWLMPYTrEq6zNcqLb4EXBOax7LgPrafhHCjvIgUsMe3mGccGGfZg
XPC8U97rhEb6lNFekhI0wp73GkPe5Xmv+dtyj73gIk09JM+usN9C1a+Aw4+FJGoZ
1gCbUiszT8lOaIoIOFfTNLH110LClvpqyGCCUbeSc9g08geRa3vRK1ch1btRnaND
4WXox055H+szp8diiHD9as6d60/QOGF8KdF+A4vpqCHzfL+skpgerA0NwPJDyutU
wsR+iYEb/92MVB8CH63Gk1LDVZ4fToa2pGHFCfq0K+A3s65XZOYmlP6MTdVx6XWj
z/TpFd5gIZ6/N6gcj9YNJjBAb0OnyT15JYDfIJnUSBiJHnqfH3utSLbiP/axMvVM
zNL4c48Tnm/iDY1GZOdxiu2Rcabs8oGHw+kjtbEyqoYqaRldrYTdqZiQDeBU13CD
3xK14O1KSix9cZmGjsHRcsmvAUdf+JNV/vK3wbC9MX+FsKyPunqleqK242IPmzbU
Y/5KRMVgLBx6Cz6wavwjjf2MeCAhCmZdV6PTvTcW9RUpKfzNjkgbwRg/PMsNUR3h
yKfMbXK5JzOM1lMM50Cwf7XGjW0Q9UHkVDgEOmG6lWSJrj95cp7wVe2RLAblMpkP
VApm9Ej0Bg61vUOtmZ6NLv8/9b0Dii02OsXurYGhkFkHdufM9RCnjkumPupqp4Fe
Fs8b6Y4WkpWn4XnHAQNgEPCzYKFKVocKneBiB1JoWL8PfDBeSiPPIPrmjxRjcEkL
ecIxsGpkgerTWqxph3DlDgOB7dsVevTNvDdsbB98FFix88/8dzw/SFHQBVzkqW5d
VGWszlaZ6QYdPhNKxrECPaJmrxbSXjJKx0yXNi4oL1JRXmXRGDS0i8aacgC6CSSt
DWhkjYmaALL1qP8B+p4CB1qB6bKF2Hk/Poz2kdK+a0zekEsj6JHxPsa/OjeHsWUl
j7aQyIhnJVoRe9C47x7MkAoeTvgkRMnw+rsFBWpTI4n87YE+CwXntHtfAViZ5pLo
74mYtq4RxF/c3iLYWA79R32U/I72YNA9l/uKiUpegvkWWTUyKAHraoIowfzQ9Iaw
6Qxo2mQ6BAWhz8ItZXb4IOGkERixo3Y21sa18TYy4R8k0IdBe8YNykG3/N/I8TPg
/4L0w5eotC3F+o2maFPLu3+/5K9YUI1xIbGEFFP9KYuv5gJ7nVk6rFiAeKE5dB9J
BqUrGe1IzWXAKiOSWgwMUWXSqG4Ibp8QdqV4T50XEZRdtqiHfSsi2i5wqx37oAG4
cPTdlWebAtT5l8KPWUSruV4GxHteMEBn0dY37JI6cYDu5aZhYgydc7kvw09zPv4o
cplB7weqwpCvzdAHFRXFkZY1EXkiQAdDN2qKajgup3GXulunz0blpVTS9z6JxeHA
GApvYLDCLf5mBnm5fsnKTxjATa/64jhrI6GBbhSZBUhDJkKXBudDpNRSeriLjV/c
+cl2D8E4p3k6X08+eq0IOqg17TZ3hVOAfHR5wVvVj8sN+8MIvW2vcvjR4SbKNMOD
C9qp47ej7SEKfF1iaDoZLtpxaBUSJnu4QzqsTYDUgWePAP+MzVoVvaQ8om7jAPo0
n5jl2Pqg8iF5hyk1u6sb7licGkq/7Ac9ukdSAkKjda+Z9M19rkgtg70ofRJVG9nn
Ur3pKva1K46sZCbIc/7Jabdxbre4IG528hXhDR4gT/dujNopUPGlDGjgnZ3iNDji
Kz3MPKlIC6/9oSSgJHgHcio9EiiHqoJGpeJEXGj4m/4t/R1Lqk4TZRQAheC7xQmf
MJ26LznBbPcK3W7ym++cbGwSVhnRG5YiFbMa2Vewae+daFP4mNbuVoi1fv3ahHYq
IIghLdKjI8D8VO7DDj8X6WH8ircTapWOmFFHX6tpWU8+pYVRLjRYtNAPSTafH7xk
ngqxzeNpeEdXjqUyvHCknepUN/U9tj3offIyOb1JXcBj2SEljZodEq1OsKOObJIY
eS3DwNc2p16hRsbJ7dH8WfYrQDyUJ/kJRUo8B1FW55XPyuxDhK9B2KNiuad5Eyfd
10VKyPSrfogM0HwrkO152BpQQeFxXZ9DGbOWQt45c22rY+e7cOGcpzbAuvOxkF3J
baG5wNSjEv2yJy73ZjmMCBbdOLZNhEg+ubNOmsRMYtso20mH2m0LmLwi6VynSdLx
IOduYcXstkRiVriSYZfXU2HYjda4OifU8fHUOERl7btjTksyPt8hxpd7lEE7PwrJ
QzH3J05877qGvO8DJxQz/2QckR0/DQ9SY73bMzpu9zE8Bx14PifLeFLaGOHXvjj2
5G4XuoyG1bansrU/OFVFuMP/BkinG9F5b1Ejuj+26DFHJSSSRVSVhP1wMd/AgzFO
aL5AkCQsX0Rxkay0Mw0tvk96wOMRmloXmARy1yH1g4HO7zaD6FGKEMQzkfYtPcZj
8rYktBw6aoiWA63tK/zBG5H95BN3HqaigQi5YSpdKCicDZUVSv6JKqJIPwRIv5V0
hU6nswQMsP0nXqp+rdgl6I0w1ZiNlOk9NC0O/Gsw0+D4CuM/+yeAJl7emK7C+rvd
pRXTLdwPnMwlyI0VL678sx99xceMzm+EwTDYriCj2ax9v+uIiaHqVz4mC4gktwy7
Yh9uU5ebZG8UOrihZB6hoBI3A95FU7TgJRuEYXJLIvIXKQPuPdIe5hw5chYqup2C
zDcRMogNx7uMwUXr5zzIx+FkVGwK7/8pfdJ5/0gsjytqLX7AopG+knRrubWjn6j9
/j7Dhr8e1f8yx0TwEb/fvuLONUxzWE8eztHPQXGim+c6QKZeJnrb7sZA9F2hpF4K
BxH/gWLigfDjxXDIn5vVFIRM/laYT2vTkFeWUl6Ot51ST5iXdnKI2f4ygby1u/Gq
lXl3w7TzTCrFEIUaKwgKQtQxw0Fsz/4jq/6mVIu3OG0+Qz23nV1+ljLdwY+lTLMG
gPBu8kYtXc7hLV6B2dE626vToKF3tO14FCgO5yE/KExth1Vn0Iz1d2luVYrmtbVU
jok+TjCmkflAZ5bsuv9XGJVs0vK07lz3CRiVpo6lHxSUi4Lk8M1LeYajO8TxARNh
T7vCGpy0SW6CLABvU9ZD+/K0bLFTRm6Hsk1+5HJwkVICbt29igwwST9qB9DnowQ2
mZ2KBQUAASQXms49ImmeHBgUEzkogwbHO3s7C5EXL88dSCh3hJxu84hzjxg81fxL
EmPPOAZBtcRhPpUYBCvyjYRvENmQ3Cox9E92Yy5U1zcZ7K2mvZuZsTKeiI8SpXYb
Iu36V6Mv2bOJ824SpZwc4yyxlYbNcD5hcd1fwYzQY4GLcdhdyWNdoyW4fuW5dQLM
wyt3SDuIK6/MSwdmH1jyFUNBa2OkC7OalFqxf31Zr91VqiwHak4v0G/HlF3F5e9P
LAdyo4fnOCnuIEYLwUvZ5n3aR0r5pK7Dh1eP+XkVkRHSZfz6BF4CNkY8aAQHReIm
bA+GM1TthbpO/xtPsOv3SUNu6v89cDBnkjt7gjX+Nz7xYbL5gc/g7unls7GfFDGK
y2gMc3nbM1yKCUuucEfd9inmkU9GvR66fdKVxDi+Z7JccP/gSgtxBI2MHC3n41Tp
OC8Db0Ve6fsHksODKO3OHYtws88fZ40ZMF4cpV9NhgR5JssnZqUOaaRnDDqo+Hyv
fHqH/QzwuMP0PJurK18TUvMenqTcQ7oUNoOy3RoxCG2EotVpVG8OLViAAHUf98fV
jMa9cTgyvMUCLwD+cgEVgDsCKm/XynSeMXLkteCib03WOKbdroRjw3F91YkJSsSn
6GmCoPv9PomAMdkr/Ge+GiRLj8quGayg4gDSZN8hM2K3ckzuKC9NBPYly6eTj1fF
sMAfJxP9YRJMol07WazjN+BnOJP5KYt2nXKWY8dCKQObWCuWoD18p876/dcSZ2h1
tnlGVUK5oHX/qMVElGlJ8eA8+MuhYPI7sUNefsqz6/m7v9nbfzb0jbuPiDxuzcyx
gRUxrgsoNn8kDokn2b+zoZweifYOO1+4yLpLrjJ2cKe0iJGOttYeoC8V3fgdDwpz
vROC4UfoszDl3s/jjkFMAvHQhYsqu7183nxRxfsL5/h3+hE4zkuZgjIW6JLDWQW4
V7LJuZmseBhDGLsydjjx5v4WYdPjzq5QkXb2xQFra2dr9DD/VuVB4CA7MgazzVK+
l4zamQt76v6CNjApx+ZKhvTs32bVKxR9D+bycdEsDjFVh0EqCWbWVsnbZBqa8FYE
lHfWyEpgvp+8zvtWA7FzPFtU1pFyoKXoPHmUK9zc3ZzOPy1PernG5I65SYd8cPvb
MJ0PgTdGBMPh6wPOBmt+JJe8OeqiPVVs96ySoK9aqPeOxrRQfZxvjpGuiNbUvipQ
CQFT+gbnS0zhCWa8fgfAiDDSM4TPNayFolxTx/uJOfYwfLo/SOnUX0MoM0T2iwT4
Dw0F4gF9L2Cdg4PJ6XsMmqVSIr4pxTwbCJGC9fDlufWstf3GSdwaqsG491z1Laao
DAQjjBg/rOovcutkYOr8aKyI9Y0+aMnZfcdsiNpHqRVw+CtznI0aty+FSuEJr0Q7
OfqlsvUA98qL3egpwrea0ILJv6089gfN3zmtdBRU62qep2teICZuDrZf4fx0Topt
ZLjzcqNyikqPghzMzvWlgFyoXFmhVuyfsoEXMBiX+4NwZJobCwNvAkWsnoRXScB0
hhEd7Z/1529niPfGMPmqTDuofW2YAnynyH2TESq3XCF4XQBQkLbIXmvBsrrSFgjV
+RnehoM8WpefCcttlTN35osfYg2uzYUM3r5CpVpPv6EdDZOa5sOMiYKv8bUgGiOE
umq/Zs9+UjZ9r0pbYNnWBj+CbVpKXx5vCqwB1BwQV8B7sdtrB2rgHY7jCwZINyL6
faX9SBU77xFjX5nHtxq9ylgcG4q+QlahsezYgSOR+aVbnxy//i9q7+yKX0snLx+J
RXJKxMz4oFxqebYxgtcbCG++ZJOzcSuoz6JJwayJddNX4wib7ow3TBZXRI2DJIb1
GTKa8JQ2d3o/VdJhVdvrlPsN3Bw1Bv0SWh18l8nrw9Eyoj8Bldo1crbx4cGEhszQ
3txqd1JG+JymISVxvGwBeKQlfbap2rB/KcfhBDpkbV2aaC/gNNLHeT4gnhV3VhmJ
8aZD0AoTHm+PGhFKc1tuNF1kILrzm8al/QLFGH6TLm8rW2KdYrVQpO1f0qks/lUd
HhYMHumusymX43KbMJYM8iIdLvV+Ah4QeBtbQgB32xFs/RhGV4SIsHTi2S/wJvjs
lLexp9CljHcyuaJ8WA0wcsvXsIptbLpaPvD5Pq4Zwn0oUzWGt0xMb2wny9tQ4dm4
zN1EXUxa5FGL+8ge6ptXgj25MZrfpghUB6+SJMd9vM8vY08wHbC64vc/vdjhvqDJ
fY/LJUhmtf14BG++xe7EvF+OAl6Z1q1vIN1Yl5gbqsiHSyo7tvc6dMSB46XELOZm
AfTkujUE6Qy7/U/A6ezZpQVkbHpv1ynQrAMUfO4LC0rx47W/W0u02TBoS7Y2Kgix
8YF8XDwL74HNGujeWV8ZS8hFDPnui60tfI3Aprmst+K1D2kZJYcaZiCpFeIqVkjX
G2f7J4+mVgx5zjv32+9Uxd9zU6JrwkiWCFemgH7i7y8dxZWryIYBEO7BYrqE0lbc
1oXnweVrT/CCJtaX1V9bQFTxC+djY2aJDj72PKb2PEqunj9+pRKp4PccthdAmZUB
hqMUD5lffVhdBsmvUc8ZVAiRPO8Xgnvh79RzO0l5s5Qmuy5I7UTORwdZcHrAUtY+
ncyOnjnHjcxZAvwWiJghnjLPo7qiZIZ+0Rklqrn5hT4L+EYKEPS/TvqnWZPqp2mD
rJgVlAJUuU+S1WhsfJ9ijwSiuPwpz2Pgu4TAfJa6Ui8xtsaI5gZxo8RsuKLf2Sul
ACMvHUQOifx3vR0S11rCR8qhmF7GlTHMOytEuYcFLyaiha9Dr864eAWiCe96A7ve
CTPpm/7iv7hESdKnWEN2hox2lhPxqwWwux940uhcO+a+LIckKMduyaNTiuZCRn2X
ugRS11KvNPnuzcqNmEiOLqZ6mvvvqjQZsxdRXQmnXIoZpT4TCM0uEoiB8LneXD7j
AvLO87IzOtVomXGat9WnUlcA5Bf2X811rm9xVK0gTyD/i14XipZnn8K60zLzLu68
Mfwdwrzk7H1JUrG9mQPFY1phPhL50kFZudqin0n9Imv9iTlUt3WZ7DyjS+bf0nk3
lICf/zNbjy6tw7OWRPDv1hzxf0TBXFEVMoinH7eNs2bCeDcoxwuqxlYhKDI6kTvW
Z4knHt57mbKFg+KbCIgx9GFuxG03KVAS2SiCHqx3s+BSsW6a2xNYsRFwYE9L8tvn
Rr3ldIj7th5cLNj3L+KODpAXLaRId8NdOmYfrGI/41xs2mT3wxqnK0CWys5DlR5T
0iso3HVTVMqmzeq7QxoutUAlzrUAxrAursgGQeDtFtXtQDd/Jfmgf4axensTTfG/
tvCBDd29aDeWVk6jtC7VKvxif/CYzf+Y1qKohgseRtwC/lDVDS66hwMlTpfdw+aM
LWruv5/a+AvY9JfglQQ0Sffrme5sr99knuHSUWd6A2dZmjofP0RyzJ8P+UJmXMj7
EIvuUxSRweO330vgPjrsCNw4+VPuTVUldOHFpcYzf9m2Hxj3uqsH7ngXxqaL6F86
FmP9oY8S9cBYEK5VQw/QRMIaAfkJtxA3pRSsIn2JbX136WUhZlzlpP8CkBtgFpUf
UHx8ofM/AFloYHjnBko+qNqfBeO+xbHlGWuMfzIh9P0gm/UPDnttlR0P6p2q6xfV
UViVyjrc41tR2MTojeuBmHOUUYOU4C6yKWazCsq1luJ1ANC42QFqtjL0aK7Mp7c5
3g8zjJEfax1ypgk0AV0+tjqxZ+wObu30TN34/F8Xcy4Bjdq5QSd0bgT1eqq1SlXj
Y09SMkTMPfhvENf+pqyqRKTNWDCYqi8HU51bOnCZlbtR0HX8EvfsmPO5zbzIYC2+
Lr3Pmchmoz+yj4PlvECOr00ZF6WypYlfQP9lWk/iXyU4zXN89vrraH/WcMF3VKmD
ZLfPp6lrM5h3znjoHZfybzA4GiYIt+yOuIzPD29mFZRbdawJNeDkgHN3rw9q30Ub
0OPgh9E7mF501Wz2iK4lb2zZSHe+KKTwBv8scFaYeOQKxQkxQn6OInxRJqnjoX3j
DY0t8q6njfyKNB3jFJzNJaIPVuHf93it+0qh2Zu/8z8ldbw8VOwMSZ9kuuSSu05f
G9I7R9fGzk3lhyO8A3ubt+b9gKPi7Tx3MOFYERmIdVN4G7IwVv5uH10RGFXwWRSa
LeiiMmRPh4OFu8uodR45PsSRGyMycw2PYNS8Fo01ZbZMNi+pkOvEQq3OSp2mCjSu
t2E26M6oeqvzulCXtPYFJWUtGJgqg8C2u9Y2oUMcBQxAPDrdgVdCRfIrJYaaDqWd
v/vgPV7fHvGwnbALIWauRn4vq1AH+LfHs04MvX/2bFe5CNLDBUFITrQqD0kvEPe3
t4S1N/U7oXsLx5ZSGCG+R2oWuQYuFmOcYoHSKAwuARQmlBXCr/xg7Ok04qhE0P90
Nh9JvnGcv/Lf5fG9Upk/SBOdiJS0f7+xSXl2iBYiYeNUxaw1FqYrDnUoLQ6egtlO
8q41jKCJZ3YlhKPxswqhm94A34kDSuw1bW8Hg4qxwae2B+HXvahJHaPGRSa1TNYN
9FElQzsuGrtM5wZPgckk9uuNOKuYane9WF/IcqsnoSlo8aVbdsTzmov0f+1a6z8o
bcXvjUqDxsuNMiGUQzE1BDenA8yfBWSB5U+tUGfcTvuhx4FZFUAoHitKkccv60NB
J8GugtJMapPYrFnFM4E1rFKEgHL/7qykpo5TQhJzWVT6T8U9ziXRKrtwWGClDgii
ROlUC5bVh3M8yPaXTIlGfBw7nAYtN9VjmnpH7J8/GLNZHOvztUnZzbV/3C+aNNTx
m8XvAyCKbzlquQY53Ul90npI6C3BiLlAqagYKEu9CLzhrLN5dyd2nEKHfghkIJfK
bMjqZ7hvQszpPc3dT1p97bH6wH6tK2gBZNJl3NJtgsUoJh9XkmlFAgXBphobkrQE
h3d+8nNqfzyb+wO68Oc1rT8J3l8TMdwDcRbaMn3thefXhKf/V8io2bDoaKPGfRnE
8BHXIxM/m3pOWAWxsYIjObawRqAvf59WH7Sddh6r8YbxkdcX2uXNsSLZfLpaduCj
amZaHxmMrMq6xmUXZp+MW7I2xNdNpGB4Q51toXpk2nVNvdz2CyuVNiPJFk9duyIW
forjYOi4Llid1A5uQKra6Qn02AnzPU886lKhJpzosNAPF/Hs53AzC5I6VLa3HA6w
OEIAKC1UnERMASH5aCeH5z2tF2FCwmp7VMZxH/hHnA86lPJraf3Ha37Wt0bLCcan
dX5SjO12hr1ep68P4/IAz5FVSapCh46M01bXM9Ba5mmeK+lTkVXt4+nh0nAYRkeA
5rXIJvsAMwq7fmA6u5byZgyisoxoeZRqLjmQPNGihlm8E/wACLQGzon2majFCLg4
syzG7/XJNyRWd56zZWI5nNq0r7FUZ6aQ7mGXLi+iPdP0+VrZGz8zPw/PKnBiNEqK
nzVOE/2wQlxEvJ9CtGrlNYPKTU96ZVFlc+0BJJeAOBRDFZGgqtshVpXNbojnfuoD
Oe5Hibwh8jgD/2aoEDnJOP4sOYaaEU+zEz8LcgCQBu6ddBynXneI3FSS04rxyC6s
2+Ny/N4rh1u2gbfJ0oxcaJQwJyiKuR7rO3PVAcvlwQi/o8JnN2iM4bHzPhkd/ntB
m1wsYqSrIvFYS++xxskpTHLISDERA5JlIJSjRGKysnS6mSTQtuM1gM5AXdbbReFn
`pragma protect end_protected

`endif // `ifndef _VF_AXI_SB_FUNC_SV_


