//----------------------------------------------------------------------
/**
 * @file vf_axi_opt_fc.sv
 * @brief Defines VF AXI optional functional coverage class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_OPT_FC_SV_
`define _VF_AXI_OPT_FC_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
msGlmB1wp7SbnFC7Xu3a6z71kmfUk338Qh8mI4HH3Mz3p3chHg9BbCE16CEE9LCl
yogYiov4N768R6Aqpl9I4OO1VwBzeQFTEDoXB8qfC530Qq4lPnpY0WQMp87jn/gJ
KQSldgfgfglWZ2wuY5VrQzhe9kzSfvx317pv8r2XtjMbmLAHq+MOX1xdU5SeyapK
DA/h29X6Q/53mI7SQyif8fSWqK4i8EK8MLmkoHmlFYbvmEpN2X6Wy1aG4C4Qk7zV
OLlVCh0q1bGHZNHjiGvQ+pwa8eOTXYzgyPn10tmUvp1gCzDFUv6iL1vlVGeTsnJP
IPFlJm2qaq77mUSDdwwcwQ==
`pragma protect data_block
vUJnUxsBpchGV5sWBqfQY488Gm6dYC2rJuj4wgCPQCTqxEVy1hbqgimeyC1volh8
skLfu+Znn145NtW5uN7cKdKYmbRnw06HR4W2JivZNKafwsJ00fD3zPfFATHSvtHp
wDxGsqnrDtPng0j+GETxwHasGYtqrvYSxDxU02ML5QAgxh8bvSkjkx7aE1Ol27zK
nqYDPYA38K1BXEimja6D5eNV8lgvQLgFIXP/Wi+Qln9a7M4esQtMXGLmXxqyp9gx
yCgGN3tig0jtAh46oCYRek3m0vi95XSs4GLWUHw9AHPeEGx+5OZwOcOXMB4E5stt
YkNItwjkTTJ/7ORbVjxe4aE8FJLXo4lAywpfFOqVLymzPd5ozfM04+nKoRbkmf9b
YchYEuFgLRBI5gIje9lBWdFFsgGJqN3DVn/8Y9PswY4VFGKzQKbuHHCWnrYf0KpM
X9x5UQJX+rCLE9iteNGbYodcCxpQdT8qBpxq3OgTh/C7BsLmt8psfDZrUXvxB3r0
Z8zbuLoXu0gTy1WI55miIgKMgBwn9O3Jma3JYon3zmQcKkZwD2DnRI90fErHDAg/
l1Fl03fy1VzraRyftMWrq22T0YHMuQdbT0qW2CRIn0/1syB7kRp6xto5zD0Ged01
tG4408qydFI6ARL9ez1uS8f+5ZicqaIlLaF1UUCFCzLQDrwMQt+qodL85lkcCH6U
ouz2SiE5uOHYeJXElKq6xpzX7yd1Tht5OuPhXBx6tywPbo7klEeZv1OjhzouA8m7
3uO8QzlAORHHK0/nDuJ9ZzgmPzankemlPa0GFxHD6WFa0l3cvx7A2yK6tWVxkOiK
V5xoNJmTG0lhuTuDq/BiZ3SCH6XRYbr0q/rqUwAu4XnSaxg3eC+6o9INx2V5I3H1
pfb6js/Xr72XQrZrXIaHAaQlT7LY7UPvsW08nfEjM/wI55XN8PNVYHP54pG31eJf
vh3xJvNxe4MuSLOrsitl7boMCNOh6ncs451GC+MzKrtwNfJYeUWyA2n0z9n+YTxg
KQOlpFKu6pLF/AXOns+AvRh8UWuvsbUUnJ1pEGOgyMf7AP5waHbQRjZpzRGE8GmK
Ica1e/eYaLL/TXEaqL6P4cB4DBrmiAbk1gUgItu8eKSG+piuGG+MRZRWJoHgj+9e
F8GAo2EUsB1Xjq3NDuGMJrr5iLJJAiDptJs7MNl2XGgfa3TrYC8GhGplpWBjKeGC
/bvpQHenTV7Mf1jhAeoJ4X0QwiSxA6jr8yVIBGSIWC6t5qRwk6glvZHbAZaEir51
mwIfvnY9W/Dm3eaJiOAf8iF42s8DARxTLNRTpR2LMdHrJSB7+ePM8WI4ibeL2BP/
336jDEBRmYQApxuE8Bq+nCbfIKkuLZEFbOWHWagdOqwQ7wYPZTHfU/4ePNmn7phG
xaX3cm2cXWdOQ6tb1rCx+UCOBovYBKoEWLyh87NBCuxdSFkvWiCfGE7mnVlpj/hI
BUQc3zz4RmcoDuD9OKdGRtIpWKgS4IkB8jGU7yA51/ztBgX09eRN62S9JdhgSvEG
ybuZhwmheZ4vrY5BOrxA5ktMUl7UMMs9IPu3KPKzk20DrFVMPKUejWSBUfY/2dND
6yy+GlJZmtJRXCBVH8znLf4QIoKksLGnSKkdPi4/SV0YnpqQ7LttM/Ky50sp3QA4
ZlCuDX8C9zVvtRJFM4BPaN/JVisHtOfJJynf31PQffjqyjVoeAGRK1KG0E8Bi4pd
rKx4qY5cA2yqv+zTQrV178ubzqSwTKy1iWwz36yALoa5FLY1RgTqnTNiki5LXuip
fZuULLzXOKzBAiSap+f5ynACjE4ujXtmjcF8zwnKp7TjJHu/k2LCuiLqxRNNOTc7
M9magJ2aMsVTzYhnIfv9qZXP61zumk76RKg1hzpNR1oWgSCDifor6AknRtN1SBhJ
PeT4XDX5ETIGJkkp+QqgkIcn8zwvtWdT7Zvky3jlGqdTh2b0z5SsU9l+d/eIAmmm
1Am2yiq7V+0ykfnhXy9QbxQjc1pzW6WgEwtca/UOvfmQqEpp5ET+Ok94t9/JXP05
R/vwwE6e3xA+ubW3I8JHhklVqlMPwL5Nw3MOSWNx0Cs82XeAJsQ9m2J6w02J24QJ
pGbKvNLEtCNGKIE7YmO8Au/aci+bjxyCvXAaOsASJz1K/CIRo/zi1+cLpQyvRahN
AeEOmfKP1AznXJmK0iM9sPwC/iuPEucSF9jeICw8Ad41bZA504eXsjI9u7SUw1CB
nGznoqOSnzhioRENe8SYlcZ4vpTZpn4HRaekx1KIftbhIk5RFtoB1NPaaLU8pNoa
yL7iGzf0JI1RVsyzNXGX7UyF2Qxkp7YLIYrJnGodKmJGc9acxFaP1mRm7ae+2FMc
jKfXyJF5d82m/ETsaWfwsenn9VVOLC0rog/i6AIm8yBPJHXBvJe6mp6zjd1nPHEw
QxJ1ctwsanPNyrMncoU3zAXTyGbAXkxp/+FjUrqrktL0BSt5DV6kOgKxkDdJ/RIt
NaFxNmBdO2mh0qd3FgE1D/1Pfk2PPHz04iDvNf03Vh1dmHrtxx4Z8+bt2srGwQrc
JX8o9XQ7tQt3ZDfoS06P/W9III0cS6r4IkE+emE123CwVAz1Mh+DLAYA3c8WxC7H
oJwpjqfN05Yy0UNYVcpAblj/BjAWrvrRqu0t8pCnueIZWkHm33Asa/4oiNKWFb7q
z9o/iJyYDx61xqF/g5GWOvmYMEET4xJkM7sRGEZICalw/HwDLgoFHxN7g8gpAF0O
rtIzmqL72MP5IQHn5Eh1YtlN21pM8zcNjUKOYrIFfYKCbawvgrImQSJmSlQtyOA3
VvRtEvrkpNrmZ718RGh0JlXA2+F5DA1vaFpcyL8gPYmPIVDL6z0ZveC5vetYhu2l
plYLEXT0zHlllih35ugrarbVzPQo3u4lXsOfiGPzQO92H1vu5+Ebw1ZB5l9PACDf
lcnstab3FZxifqMaQqrh16/Bxfqs2ZmZP5Dnc53eNy5tsrueFhAHPJsi4ckSdEio
jAoULxVLVUnlKk+D8dGp3fDtkPEw+fijjPjGgXUywOmzLAW1g1VdkscytdKCw2Hr
atKIvq/kCpKS+7mjz2d+XVaSJWa71ZHQx4SVoeK9StXDJSZPYf+6AShNZQf8TNFM
2t+p36i1RoF/SJxVZi6sKdPG0/Mwsp3VvX+KcoqRxHGf21anCUzp7ys2sZ0c9rOH
KsnsF7vXBwZyG7NmbmDA54ZrAdtg19+EiIX5Bzkq4FKBugt85Yw7MvAa4NEZU5y4
Bbsu0jWahuZlCe44L1laaIXSZBRPn9DLL02KyApY95+L/Impwdb4NUOpeQmf0tZp
Vt6qdsH85WX21mScGEuwLnAqJ/fSneCI4WehzfJ5LubTdSHgpiLZGQDuuttykrv0
8WuMzMtys+G0HU/b1pT96jHm4By5NAiuB7Ki0Zz+0VMkgPvxMubAjsEJ90pIGQum
pWwBbXjfiscGhEGrx6r0T+OLQRAi6Iel3xtW0rAFfOM1xZ6+Plp8HkpNykg0euek
OKj2+F0UfJCMx6z7n5IXtIXns9jggEiv8sNgU4Ytj5Su2g0YzvmijagXNuMkbrZr
fUAtWABtnVQNQkQAXKarq2NSByiCc4Se5h7n9YcrTnq8+aMENDdyKnmAcdWz7t65
CjMpWgHgUW87AoCVVBtDHcQ4OmomDQ+B16y0IGaIqfT9f4MwvJnGIrzddKfd1Zgb
KkPSaQTygks+QDt2Rgswl8VJ90HCtDeRgW7C6iZPygaMZNnZmMKisZErlFEf63oT
GNNFa9aFqYjfEFxYjzlzW4sVRLD8jaXiofUApDAedsEM+Ic+/MMK5EYp2LJjUpy1
H3YanG0jxOK4sH3dZ8OjNfrSxXJZI5yc5MgWBSEvQigf0jR9KWw5KRELvnCtrSI3
ZHQx8NOtXxUprf5uLnWH0/npXCQUibwg++R3T/mtScPIBpUBQrkfXA3rQtNt/Riw
OXjBKy15LgmYrOGlD6RiuNuL8iVL0ebXngX8p3DvPsYAdXMLjEvyRxqBQWMMxq5J
u/Bye6cmEe3Dp/FOFQKdG6g5UqsbGlMcXXCm9nJ84Mya5gLlnYUhFw+Q+irtOZLu
LRR/1tSN8eKePnN9YIZv6hp/ann740Xf2BeViva/xvezaSzqb1TRScfi2DvFXNs+
jUjR4eNGVRrLVJxpFCEw0CQ/RpdM3dRMtY+G22kyOyg/T09O+Xvu+t6ifJaySlFO
PU2OgmyUIZPZrUtam826EY2K6P+B+SoxV4bI7vOSNyYujuNUM7qixHKw4yGwLRdv
TRr6PwKhNut2QUysTB9K0DaEKmnlcHNClDpUldBIDP4PyxBmzECIW6r+igw0thy/
ROgnZiZkZt85A/IggRR2IhSaHPJqJSyVVXL4Vr3BmleXl5+l4H5mGvHwUV70IGIm
R11S6kkYFd0PoXiXhWArONjxVM6CQz8vK9U+qEDE+Z+LZLNADl0oh78qgf8c18N3
FWg5Yt76Zasl0FkJFFg5kJ4rpcpQP7e6VZcf074UPwxyKmlZkwTc1M5NX6lOqHZ+
jAe7DOPB/vGdyc6kTgQL4uqyeO/k9OkM30i01bN385MYZ4xa1kXZfe75VYT24boP
KFAwB0CgGifdHWz2RO81Up37yKBzahS5Uu5TsuZT6o78hxBmvLaowZEV+kUt9HC6
7ujChVoRkjUTedPVEHK/14HBb/oZzGyz+UaEQocaUi2Fg12rC9oxF7WCBzy903Qd
rLBS8gqR6EOpNodHpeCGPBroJgT2AlI2Rj42x1J80UROLU8Sex/jcEg2X+Pq9Yyx
gK9Xno/Mb1mVXMGAl1tAylOdkrBWkyK9yGgEXgj4dK4oZ79JoMLupZEwHlUAuIAU
A4mGsm6+rYtOyVYi8WKfl/bCrLhr18iXVjOIo+TmBuXZY73i+cqY6h98cwAdxQc5
kP6Dv6P2o2JmN/eQjrrgkndLTCPBTm6fC0XU7iJ+AhlB/JX4XZc9eMqbCfQOgNPJ
jKgGZre8HlN8AmTrUan3rL6Xe3Cod5MD7xBGPDEh32s/2/trqnsLf/9flAJbaEzc
pcVkqdOK1TsQS5AYECkgeA09F1xilQPeHdF0pgnu5akLJpoRs9QO3S1eja9qkcJZ
PD7AqMUXnSnMBcPpgv2uVCgbPRBlGs5pmmKLy0Yz8PAAvqEUZr7//zhIO56Ai8oN
7EWheU3YLFy52FnIPlnlvlOokQJ1J0SD8haAHP+oFLpRHRP/NICx2Ae/X5zNqCXC
dZIW7qjfqzOiyZsG/wtZCbgF1GCnCk4BEmfyu/b0/Hf0H9L2F5TlVW0ZPQ8+rua+
HLJScR+YqCaXEQDgF3D3eiJg6RMA82DNnBA3oOnxeVTyFK81nUuOqPejX4d8+zt4
sSzKW7TMnn9Nyo1E0yU8rUBZ4B5kBQyEmKQ6B+GDJkhscURy3SZ9Qo3WvEy6PBfu
V47Sf/PQEADftOYkNgMbEJaDrVCJLGi7kmkr8Or1dlBDp/jVTDL0O1ZLHhCrtv5R
AiGu3AxZCOPOwQOeN5S4ehXHJuVNh8SWx+EZmFhDafLmuNUXRpR1bdUFgEdPARlj
C8XWS6e+nWE+ASEg8K+o73sAkDyiScRj2BNOByYCgEBMJDenqJixpLtzS8qO/Nun
hvzD3X8Lb022azdccph2D6LgQUFDlaSKjQeBEJ2T3eP1UD7aiJuWmOgW5+npFb4J
KP8vzGY4YNbcgQhimsVgL2GwbYJ/Z7mtzSDSoyqXVNeP0WpRjSwi8hIyfBr0NsgF
7M9j7YH/va3lJTWSA5PR3allTGj8BkOGxxOhMUmWbeFFagUDHPYzDRWPG0NIcmGm
B/pJ9OTWkG3lBu8kXjIThkfoGXUaB5jHG+MUIanNU8Xg8zVJpNDD5SW4mPrC0CyC
i6/MzQN3HDKPXF+RJWGiAuALQ86uK77tnqHoWX6NKHdkPw0YDJG+wfWwTe9LIYS6
YJ6o9yvQY7cdtprqRlsQmKpoerj/zPkbTmQ12Ux26MdnVlGDjJq1bviXj9PnIZLj
d3Lk7zr4sMjc2IBYk+NbWl0lE0IugQ9ZG/9FVH1D+t4tyKQH9x0Hywr5kVAmLMmb
9Uo24/q6SiQATQXydkvmQqlzma925eslE0F/WEYm0NIyk0r8pMxvsHWNnEALH4RE
2hYbYU32LlRs3T5BggL3baoAruptKlc2vaQegsZ+DgcLD80xyrXMEeABtWRye9Yt
SNHSZng5yedNHOi2pyu+uJzByZ4gukzr6FX0/UWyixdlo0i5eoJtwRqKyRLdwxGI
ao3cNQ5y+/nQa7gnm4fl62OMWrO3DOKc7pi8R6hIJE+kvG6tAkfGs8zKKFeHOIIZ
kMBIB9Ca9+UDY7sgL3URPcy4DqyX7wC33bubsaAiHvJWQxEh0SP21CKOOtcl2vPP
EmqmSykF4I+/xtIMzlnLGrxDfiahlXwds5hP2RcngIZsCjBwK78TA9m9P51bK0AF
wb4lX+61EagWlrvaqmjocEsG9fcMYkvMUn0KTDPSY6ZhJJ4S8/lJARoF3OGcqqOJ
XTmJZbeik89QJ5HHnYfyyTnStV0o3ysu3bmSFUPDvQJ5yCcVv3T7TgPrUcCU0tsi
ybfXrGGJx7dYeoBV98mpTxmkKd0HuN0ZN+GAFsn8sL6zVZknGaRX+uGFiWZQ36y9
VOvak9D0FnZMUZ563Jyj3Tm5IlUDcZrCabkgx623z01opSJagqcW2x73s3kwJVJb
OX09OPkwc/hLYcLK/zFD4vgTg0rSRTEF0gNUSecOtxom+BhRbQorM5WCK7s6pcar
zYMX6bUGJjwO8Q4XEpKitE2UTLGqWF7f6nkLX1cAnTphcGYchkct+NUp/gn8r+UH
/5JTMFB5hnCEzMA9vnyfe6mhEMC8RTc1To1OCgnpisxQHx7PGn737VzUf5uTMSIg
E36aDApewkvoaxsKhHt4MJ6Gb6jZQ1mHDT7x8Ir3mVA7++gKosBG/dZ7b8n5gU1S
svkTOV+fpr0wcFqaIdglhtPT9/FgVMBMGQbU3RjyRcvkT8nkgWkzHQK+dg3esu8h
We/rHf4+2r3wPAbmZqu0Zjx/Lrkj5E7V7gPlebQz0DSxNXnQs7gygWgq6RHZ+eaN
u9LJZg57WpZgMHIUsYvdzd/plGG/SuuEDuxaBCqDODBPUzzCJg/yq1C6UAZ2ICza
hTu/b5T9B2InUmleYIGFhq4UtG6zywQJmNOJ41tMC3npxXam2+05PUorEGETM+O1
bUIMBUaknWR4BnT3ABslStUqlew9mb0I1IeLqzDksgNhDbjiwGVnNCJ81GO2E4Xx
yvpNXatRYqoXHky3f3UqBYlraMa9PCdRSCGw3P1FQq0GsKLM5mLPqlNJ0/objpZr
LbAhI08BMuUQTteXBFY687t8x8khU5sBSrNwiInu0BTqkVjWbGCY1eLhs18V851f
shFB7p3v3GIE3eknCgt02G77qILFjpfu15xjCS7RdQ+KargpRPNKAq0ggswSp0td
D22MbhHKzQ8c3GVOaQ+Uiq/jDRPpPZQllkrV/UZLKNpKH/jH1jDPXmqIais5RONb
cqbckw0MVuZqgHI24rnON9C964FHZMuOEH1MLTieV3/zeexCcntNJ5NLcivKVX3T
7+zqoiEp2c5Iu986D6X+TK/3p8ZmShUBgAF8qQlrTgpJ2uNqSEObsdq54wWU3JlB
GnVl9M7Z490DI040HUtKJBqaGvWHBhV2z1drvvk4w4YCAT/ARKRdg4VL3QduZ8Ds
csWYR3VlVTIAQowv0hrbUkB9vcxbznZCWbDaC0KMb8RHUBpcwMgd74nipd8CDqEG
rsZhxseqd7YUAphX3EBGvx7W3ehIhRLWZLPyXLE4mdd12kaqsNZGkcVAtb4uoe7A
QLoQ+cXIygu3WNzMZS7ASOdbrSCG9dI0jx7NvVp4tDaoZAKX+Fsrvg+2T1yMnyre
YWLL827zfhyqqjtPFzgd5s/9F+FhWK8AScf3y09gPJHZ+5kFx1y3LUzTDaswGbJz
d0NmXl5aZzpDP7SP2SsV5H+0nsKMhehFHFXrt1zPrNhLDInCOOo0jOB9DFjMmsch
dWzYWVC2W+vXGlGbi4rGt+y5ImDUYsNKPVBNsM30opHJsfXOOZYsGPyK4GiVUzby
nSv0OhwAbIx+9WZ1g/yz2mp0d0MoBDMPj01ytG3hjklaKcFoOUW5qaWdjG42U2mi
uUu/fiDM9YsnUkehJc2C9YJs/7AgTyG8i7H1ljv+5FGQOJ8juuKWRAXmiCkkLlVj
AL5rZeGfn8sU9sSkeg1JOP+hUA5mHlmii/IMupLaApYT0pqGvtxUCg+5zk3XJGx2
6NWpRzK6qlQ66MI26KBap8jpEo76HREt3MNDXTVk7G4nm1eGt1hBScgE7yok7xEn
bz02oqbwFXTpb37uzlMPngPdNGAWA4qcl1E8a047GsQo90QMLvLhkqKt3v1AbIsc
EN7CKnMByytT7/uDJDZQVlWNlR1HjyRf+QI8y/pac8DZcAq4j9fhdwSKHEFMpiEv
QHt6WQLJGYizz8NErh0cXCQKuPBBbv+rU/IDo29iwT0jtHi4NPZF8wfU7SvDK3H6
64gj8BdwpNSIDDzYpTpJVfI4zhSX8AB2ebhzJ6XSM3z/7z3yJlXEpP7sJcMfE0yd
Qd+/20SnC7f4fJMyJq2nup57HQUg6gXAeAwBM5REZ8iuqRzSVBdEJLV551zmJjc0
YJXLTd+H38sdAa1X0SoB0pMSjyKhwGaDj9qysMtABPqAWXEPu4Z8Tpf/b0GQGM0O
kZ6YbXjtjvr7J7yqpnPK1u/FoFGrJpC/JZ1hGdoarrETbyN9nKlDJWBoJLxbYGNA
rN9d88m62yRKLAsF8ATd5mbWlw3DUyzGhrUSe4X7OFPN/4KR2MpRLBI1XBSO0Vs/
Au/XpsLwpyQ7J3fD/LaQcye2D92Z7hsXmirtaZ5FxhPvqWOP3/m7n8jLoAtRkCte
8DGWVJkCyicPzhdTiz2U3WIXFAXxJdZp+vFzHB/cTIUyDkAHdQsm2/rjNJtkhMAe
Q1WKYDFVHFn+UKPFQesCjvvr31ASo8WbfqV1OnvX6c6C+1MVEc334jpbPnpEgul2
0qs2MsAvEJzpi7hiSw+dfvDdamRkwVi0r19UaYxKNhszXd49fAcrj1/nyCNcLzDe
K+ZSQ7Iky1Y6UcnRX/9yjUkZDXLvr0KRp8qFnJU71JOiQ2vKAjHxlYUnC8gnLy+o
pAGqtTe/OM/Up/XKFNvt394bacaps2CSeeW9hTCy473q4xPElRtmy85eUzh2sp2+
n3ZDjS2EqZp42lo8wMm+69p/Zddo0Hlsyx9T8SXC0ofmciwOu/16tE/fUW7lyrwI
G3FHdIC6RVu5DHFfK/Ze4VfWsCCH1fadolx5/rSzkRs5UHCpCz4ZNzDUs8lTol5b
hRooP1TruZ1gxvOH3qLGiirYAx8z9AUkZKHEoaSU3WNI6uY40ayc2qdAPL0idhUq
PcB4/+1jJ9Wpa1Ezm8ONkjkPp27vH1LAzUImrUc2Zmj2IR90nKSasz1iV2XirYEA
jqu6udQVElzCwrQcxxAhp29YITFeUBZfjg4KHFDdjsH17gpuv/V352HWyqXDHa/p
Qf+qIgLPcRaJIDLQyRh82q03JVsb9dvhn9NtmQqEv/0K8nIwZ1iDQQfNMVWvBo1/
nIufcQ9rMAEF2wnwcARh5c2st65PuD4nAM5i9QYsuaicctqnuFXdvnxaXWftgtG+
ucxXCzilEZiykgJMkWTP/I+QqG+odC5fajUpFM6YFibnbOjCmeYr4M+IxtmcuJr3
TEcCnKm6iUSlzHNhYlNa+npGYlc9oHXM4sswXvQbgl7DI8w77npQ2h9MF8VmYF70
crSPSESd+Q/M5+uJIsGVYEw86PxJDY13Jt/ZRjKP0dENgeM9Lt05/Sqivn7KBgC5
f0nb3BcIflhwGdcyueCLNFtIu/x4HVKg4w++3LIPCWI5jGd6uTAUgu0Ys/fsv+IE
9P6HFKYFN00pDHtn3dObxPkC/tc5QcE7VkCfOZ1+edQzmB9/ztl5afRamGMGg1Uo
pNtr8TnwVedYdHKTDS5hKIvjhRYLgLwx5Gr6SRwEv5ytBhZsIt/B+Liei25lhRsl
dFeoGdbv1Z3y06D6QvlKtsFFBHaZcPShsGwyaJ6nsbXVhMWyHNKEKsuw/AFhCWyT
1XIyD9aIEpX1KY4Hcvti9ZiOTmz7clrhsQAK6esQ57iqwk8YhLJXE6e8Ja9uvB3h
egDAGXWIIta5BbemDrV809pVHAAcScSMshly8wLYPS6TuWX9WRqYbVQEgd/ZAJtg
uprIb5I049wwlprRDBk2wkyORbuv+TmML3Gv1fe9hGdk+cgXLFrQNOT5kSyabr9F
ebew/LXVdbMSvnFq3Ip8psO/IHlmECuUkpKmS0TIQE9lkZlxU/Ilz2S0rrb8jiTx
f7Oa5Zdpq97xhAxWN1RUXBkgfdJU7OCcONyjT2Jam4N6YvTcyF9S+Cv5YFKWhwnn
qBZGCdSx4dLRYlKOXGMvOeFA/nnRlJPEDTrpAi6lJWBpnVDPCfn6W3H1uMCfn10j
6UogbylbpdVALj1+MgrVZ7+1JMGiqIFAqbc/yWdEylGvIdPp7yhIPKOqbMYY3Nk2
IXWac0AZuN6bPFPL85VzGNfxC8G2iVbcdg0/1DwKVeg50ZvMNeFp2aeoOHToo3MO
YdFdpd0tzp3cxGK/m/A3JyZCpnAHZbQEYXdhBm47bd5kjdwUyYCKcTP0PJHJwzVu
FDPmu2Gp1usRUejtTbbuujXdkFX3mQ8DQ1LtbxYrWNhV9aJCbTOjnpvgTwcuczCc
vAccrILC2r5ceahsnTUi/VysUyQCZraJTlNv3LSvozoDOONTQga8N3CArfNpVuQn
nlbMdeMrU++uGG1p9mgdVkQtGCV3WEGnpUd5fdxhdHInr2BuIygj0DghgkyvA0ff
o+baGSE6kDC/YXYTiCPmMhhMadj5BOr17kLQBr5evEbIEe8leMbjVgyfIlWZoaq/
F/HOxKU4p97pNSHZbFhKe/ZlI1jGBX/XufQHjwEd0ZvOmEoqxBhL3sLw1fHX5YPA
NTdbREU9J6+9+f35nvCPGsqT7jhh5Cz+rYmULdHDbBEuzAPuPC7/7pml0F0/vDis
veBToXUPw98koNZXigUSSvMrFNow0kois54VPW9vGlFpzcGhSPAo3DXwM7AmmU/o
yUPkcqFU7+qc2FviLoDOFrLl0ywOLGqr2cYMzzGoHOO2a+IbSBrRzofsRyUzrf9n
YRhOn0RL3O138H3wT8azr9WKiHgI4IICf7SnjjVNEeQrjRObyV4wY/oc7jfxIHyb
STEWdarVQugABNDku7G5wwpewFRc8WGe2k2w63Fek2yw6RQvK9QQrjK/Q+t+3G2F
gM00lmdtqhy3R1Y4KbBphbMrScJzfBeOBlcP1pNYR1cCLm/pCiHY3pUYl6/TxE0n
LerrgeKH64zn9wCTEpWFAPxo1aSAxtV9qkYYIKuy1pAT3yEVFgXGv1d5UjW84qnR
08QSADgYYgnsoQ9RjhsCLsjekohPA1beHMe+wYFklApGjlqY8dsJXsvQx4aFChAh
LtwIMYaV/MGHcAyb7VDVJyWP2HQ9nu3cRr38XGu/PsKAJ5/J6a+AheoNfgcJGQSg
cJX76kkAoSbgpsDCi6IIi3Hz24+8RpELcZ6teAWTHtVFy9+3mvxhLgM+gPZNnqy7
e7zo7+G6OVxl3SVrNbPoDnhBwFsk96jas/CT7kXnLH6tG0jrlQ7UBx1cIXCyCn5m
/aY8ZEufxkdBP7VmWSy0dfBSVeokQf3wbd6WMFHL9YK+XUjI//e4FAN1lrBTThgM
AlhZdklzwk5DEuoiKXWPDP941K7LV+5uQG8yiDpQqcos3TZGnzV5pvE2k3VwUH6d
7i3DbgxUhasA2JR/BV1QpfWTiuhH+5j2i+LSS80VrHIH1WFbjtey07SXbV2a/Cd8
thZ7gnmsb1ecBAls7iGGi1vNU37D1QT3cWXlOFSl1T4b0/tMgdNcaRmd7iKpAJjY
JYOCycyO2MI9RaPYPK+PBE8a78pSH3f59RHE0cd/oE0yytvM+iK/AY0AQBoq8Nhs
wPbshyCWK69Iv6mMCu24sxZSMzk+/TlPUKF8UeU+fz9+ZYYv25kcFJmK+R3cyzQ8
7N7eGboU/UTkUiPVK/E76jkwMh4fyR145ukEqU+3fyeXziMt3o/ih0+hDL+hJIcU
o5i2zTiza2UlZQXH9AuwKfp1m94S6y/gSg1J0gyUIog+97GNs4BtoIJY6BCoUp7r
VhJ+LqH+nRjY8Bb6lkRydAerxhkdOplIdd5eaW5c15cdstABGh/G7tWLy1geULjz
8DRaDIpES9gkz1sugGsUPb+CUG1gkd8K4vcHzzVuE4ZLqn8MwaW3hpIbq8nZAaLi
9SHXNyT5MQo7M2Se0DoofCga6BSynbvEap3nV4sHnTGCSMBtkV8wSbv0Uglw4H8C
2sDr8GMQnxgI0vTUx4x2EH0iP30p6M7NT/Nyv/Xf1Zsl6JsPTmXm7A0QL54Q+s2P
fsIIcev8H80Nmr2SgRbi6Qk9IRjghL6xwlQg5qs3Ew2lgxTBrPBrB1GLJuiNzUxQ
6nN01tuJJWsRfhw/nVOJWwdkrdFAQAV8D1fCme3V2TE8i/tKDNhU9zAmdbm0sG8C
d9OEzfhYBUsXP6cZIXuZ4lMW11O2C8BHvoIYo0d+AikpKHKZBEWO++SEbTt1MiyW
s4A67SEUmCNSBk1odTYCcCAwRP7cKIzmcPiRGr7lqTrqadckY5cmyjDiHGxJRpyu
oQazxgaX/zAop+7Cs+7Zl6PUSaM2K5Kyae72c2TRHPIfXL9L5xSIYsNPC1go3iG7
54al7tE6yAVj/xxaOvAve2RlSvnVrIr1PXK2rpjhwYYCQtnTOSykMUbVP0LN+e5k
EecKKnBPcqnCirb6Yh8EejZmHz/9+B5H74qSu+5/60cjjGuZ6tyG/WeD/nTWhnrg
qVMjZrhO2Q6dWrOF5sybFWrqHVacdWHZLAiHz4HvJFFg1HOt5FJyBArdPUuc5Zax
hLlSIH/dhbFgH2RfYH4HKpn8jmCYLGlKo/Kk8Vfi7mPdGFY/OhBQPW0yb5uXEgW5
raN2j1sD0eQ68cItnp8DwpNgdQYJhqEBSKT8melZcMU/3cPH8ekeuJ2rorO2fQdY
YMOMgePYFnJHhkH+CTkPoayRSpHn7+h2XSUNlIIXfBbUPsHnMcsAOyYzcXXTnPmX
qK9t5eZWKR3844avVfn+OZluaItdMU2PNBAahnp8yrh7fchawh4a/QBxUYw8NYOe
ke4PrHrDzBJRJEnzOaTOgJSyX0o869TZUSAiRenahfKytMI/wcB5BIz/8ge9i2ak
+LY0MvjmmOiH52uZ6pdtV9HZSUg1YwQSF1Ko40eTvb22xrc1MhL+h2AQICn5r+gJ
h8gvbhpWn7KLtUHXcSnQkMmr2PU2HK0NHQNBF8Hq4Gg3sQVPiIuYjKF8Zn/X1w2z
1htwsYMyc/jSlQlwoliL8nHAJE/v3MTNQt9i9z0Dy75cA5Qz9NnSX9o89NUoS+wS
JhY0C0+pJO/5CvqCbfyIpxFZdzr1TLYCZnHKGLOyxSARQ/TO3hfQbowc7aZNkoGO
Yj+1OjIqU5ikB3BXMwWqFW+cFy4ll9yPcSaAuqePn0V0kd3RhMeZmsu5wGsh4rhH
2U8pnvNjkFfLtPP1C3wbZ71ab/HhPZAyh7n5FX+jWBwJ0+cDqwQV0+wVzMdhJbAu
c2slH9xeO0fnnNcnGGf5VpQprNxc410ztkGYYCjYrdvwVoNqSI9BKsO/BJUj2KPu
fNf09qopck2WNA63Bepwx9bqM+tKdT8pNBVsjPqVx81EbzCmUivuaLvQ/Lp1eIRK
U2k/Q15yJPhgFgulTk9j3I9E67KIBh4hhG+dhY4hnTws6wls87AR8zszkumU4JUe
Gk8qCm+V1VY14zx0sjICTHa9FvtDVqW5mHxI1LNMrGxu5fyGJfwSTxObu2v8EF+a
hWRv6TwyPZYwY1N/w/vG3a9VxBY04VuGPkXhrjXi62DCioRk3KlCec+XFdhGc5eM
r59njRoU09B9/IfkCULIMs3HzmliD/Gqsatg14BzdJN33iHHfY6TqF4uWGeJs9hK
3FOF3xJxkCC1nIB1V2HfxJ93TDc/mrfgBK/nQ212nMbQF77g86KKGv1Q6oaSTNd5
orzfm1lsr2uLfiarV2nopHkFThml699jOGXVbYLRDZqGyldpIEEkockWO8KQZIrb
nGjbWRItyX2PlLUgJ0Au/7DsaR22osqwYRSLiYTh+C75MEcyNOkA0JiJk9rBcKec
pRF4TC1ogK8VfzSncom87cUUyolB/FzeSsoavYLAfLJld5vIgV2qJXv1dGAETj0M
y1rbHweWwcido3utXdRAdIhotCbe+ELno3//hqmuAMMvyzcRf7O/OCqmd9Ywxnk/
D9I1QH90E2XwJeXZ63qoxRrtX1BlJZDMw9tLQnIRcrANGonZNJ0c/fLYT4Y6cVeF
Wguw7Jc5sleTNqylvyiRGVzy1Ewk6Cx6f0U6xD+kyhVrGD/NC7Vl/WR6D2egIUN8
06OhfBcCta4trTIsY4MZkWR3u2eR1jQTeWiGsiNjj6udNJ9YXDWR3sVd22OFFhrP
OJAdGg/yPQ+W1fd/r6o8OhFXE7hrnScnuZzG+TTCR+uURNYQLKAnCdyxvSbCaH3I
SP4V5OL87Km7ynJub7aomFlN6GD2e/QRETD0kpzNp2rCDJPV/ucwdTFXh7CBYQVG
FVf1I43aQnCVrmkJ9PKOMhCGYzoSXH/H0QLxD0hO+o5Dm93MR0mijJ6bvHt5Tn6l
LqXqRu/FOoBAXrdcuvA8me22mmZdZDMA8YqAB+fgHw2+xg1J0ICmcvecLiA7kUlb
Rl9bD7caWa/ysKplT+KpQ40Uqqruv6yOlxAhcYk1W798aNoz+711ej7LP2nnW422
gJAekDCFEmmK3Dp3glmzZFdq3KNzEwtY+RqbSSv8iqVoaofqTPm1da+IsgKFqcot
Qx6CRGCeGjhsZAyNPJSFg3RmmwTUEE+FDwnv71K2MSbwIIqg9sZFwXhf1eA2ZOQ4
AHEjdPJigvrCUin5vLJnRmR3bbqt2+1VYToQVfknmvewliVQXvmhltO9RUik16Nf
umuHgOXJ25QmPNgHJ1nHUBrIP4RdL/EwyMAXlVlmctYfxfg64YB6gJOt/dtVeUMd
w6NJbquGJV1fQXbnoBwlMI7I1rAnk0z3uAhYH0C1yl+8R8oNPvC81T3kKYN+8AG5
o4rb0aQ4ELk7scf3LUVJypl0gGwd/IDPzQWB5cJvBcehO9GpJ/R9R/MGdrLg4vHo
hacKxCVpEm54ResWYMS4Oxq32FpsAY6gwF0d2xRlu4uGbdnOlplWMKo7vBPETcnn
7A33q7vnZvpCpY+MuCYKcalNG36p/QbxZ2J99NHx/2dlw0i0U1nDNMJVW006dHU2
Kpi6Tb5HoI7OvMnDmMa1wQUw0qscPsfiQhqaWmeMmf6B2XUAkGVtfV6h6+JcjS0n
s5gKh4ly2MVS/7rwwLtmu+uIYM1QvYfEIn7fAsesnERPlfpda03xLGP8AwOP9eu5
95OLeU6xuyXbRWrnsL5YyT2ty7vwzmGKqVvgYnej9e4fBXKLeK9bWFZCzeXRJdmg
bm8XLFQ4xzE5AK8QN0yMeFQs694Cqik3Hh+hFwkHxFys/ZSLakszsasXXEQlVuDz
d+LzvBgkatV9NPkS0g4Y05Tj636qfgE9PnYdR2vu3FenH6AnJlWGIwRMP5XStq2P
VJYG7l7fobvGYuJ4TN456EeHggDiujVxXLq30qn7QgFE4MV+8r8cyONbOUBuVHzr
iacCEuoWsHHvhunNLKOmkrRTo0c80ORSs8JJxqffcARg97PWKcG65doD1zRV8ZJk
uK5pKQcViyY6ZQU7zB//labjPX8xAooL+XIqDLpfaFiGbeHYhtvWg6sC4L0q2zTm
upivy90zZs8pyUahmZrGUj+ZsKTqVUaTwBtTRVVz16SRz740K+NSBh6csEoC06UB
PhL9/gEnTaUazFjyvpWEoOvWIDAbUQxrXpmaGK2DIROxqZYYlzdC0loRqcSNkXXB
3bHQkvOEA0VdNCMF3JsTVqEKzDgxeb2MHU3bLXo8c462fLu1jmdBcdAn6gSs2Pf2
1zUhtR7dBhYHh05JmK0Qi2iVgrkm1bHXEgwU26SwWkI/r4mQqUgjzjlyigm4XzeY
jQ+lIPtcrIfBtHwLZeqflRkzL5M8JTLGg8/cYyoD839LOnsOBEkPVL3I8wa3z8d1
uAXOkBye49JPM11kT9zw0X/RZYmnGT+gZA1lSxR5s5hkhQGPwjSvah+W9Hu23U6a
gXVXNsp0Lp8LrSFgteua3f4ywJf3jJYFa7SWx9rSge9qVcUsVCLD5fyVCFJlSSjF
d0og8osBgnZfM58hCMPMkh46p5tT8zMi42Ff+IdOB9R8r6WF4MnpeRtjNMfbcEoX
VT5d6z0s8naCH9S4Y8YKXcfDnq9W8YBtGTPZKqVEBo66MOePc05SfZ60ibVbwg+B
kIEcARMbbtpU23CplQjJcpMclA7AeHxmjMekkxhLQUvT95pxEhm19Lv+taeUjujY
7X7cgKymUN+WhW+kOopEcaKhu7Nh2p6QbHbaqGSnXAlNcuipRBHl8vSu3ZFq7WA+
kW0n0rKwrGrIJacgUh4OinTDddSIMFN5fah6/oZx8XrLcDIdC3925B6wIzkkFcxz
cbVx4tKN32Ju6ansRVwuxl1Uj5T805RJlcBFm2RISId8P77M45H45KGaCX37KyHS
VSngH+EhyUq0Cu6+ehIMK5vw3xx1f0P+MYxOtFXhzHelXkflchmqVO9gBpfgsU9B
/sdqu1/VcMOFzTj0FGm3GzPzj/bIVAxNxfw1An7RLG5yp5sp5Qz/lRoynW9UJLXO
1g3NZkiLgBTvsWj8jcxuao/PTgtYIB3U84FldcKJBYokpz8/5Q+dKvsIdTpuerij
KpElEsmoHihcDHupBTeOA2tS15c2/WjrnpXVXFm01oFAF8BwkZ9v3r9BQFS6nAJH
ILSsHipeIvMV6EInyxcpWQhBAGYfluQbT0MJIi9Auv0syyZGeRHdBSDmuGTBJIBz
us+V+iRblpm1mh24RDZaP6Nm4E9DdQviuPmDHXGHNHOVxuttoMLzurNhbgCWWEgH
2ZjH5U6/WnWLo0hGfwWUv6/hVWbmOjo0YGfQfcbn3dKP/yicOpfi4yHMYcqeU4xx
6jqtcEj2FFik/EV4GQurLwegyjIkXUcTT/xdrerj2tg2VrYqbQPTW9s9PE1j7JEI
TmWhtokm5fETAl5bSdN56MFT55j7E6vKkUfxgPRqGFtZXt2jrn2Ln+e5KJaVBlag
Rl5oq3m6LkN5Fnmd7mphGtV7u1xXheKy5xCC4x097PNw7TNX6SFlO61tBYFy/v2g
brmsLRY6sERb7h1idFRcMDfzaLxYfrfH1WrmSxmXf8p2z3wnb9Q6CUD+g7oWXgmQ
/4/08ybGttL8IhCUFqAt4SzI60KXR52DwW1Twhk04Ibs0JZu6H6vD/zz76Cu8CQW
yMeIwmbepmoc1bCSSseIWLPiLJinA1+EIGMnIDfJ3hZu77YZib42Prbn30kwjJuW
YK8TASalUBkYxYz1hun+qrFu98PAW16JaytckZ58cDx0QjJDd4rr2Nb2nrZToApI
Sp1WHVWfuNAfptEY5I/0xnzyjeSx45aa8vkU4yqPa6ionHlOsLp7rk3R3t9wAGZK
mVt2O5tHbRFMB8CE80jty7UllTGkjmy51VZoSmBAm+Gmm6iA/frU1bTMqCsOagOi
uxAL0VcShnnqFgrMSeWrfmb3DfLGUNVFlrtIWczoAGok//71KIhHvqX3zr3SJcux
Nl5LbiFDJpTaM+8XEhcVHLMjfCSBPL63QJ1Kcvi6+2BvD0gBFdKtHzeuJJddjfpJ
O9qxDqb5wPyOD/tPGlVhWzFCAhv1mXrF3zLLCChohJMCYHw9Xq5K7zavRBum4Yu2
hjxwi8ivd41L7u6WcqhIfrCBgWB08J4iMlHCa4Xi5erNF3SKc5sFZrtb5Qrha+Ny
XeOcklwf97teKj4Wd0FK/CymdKUKBH/gtu+7LXInuh/2ROWHRCI/VsyEL7yXyl9S
s5yiJ5SeZZUsRfIPyj9IwSrMXz/VZaNSqbUGoFDUIMBG0sWVm1jDmNEsPB/W0A9Q
p+l37L6obiKewC15dh4rzSs5uxymJWnpfW0Y9ZsJbMWYyJFaAL/n0XjY4QmUuI60
HbNx4uKO9hnAZ7/7HVPT9fJMvEPxrf4/2RP3MHPzSmjBZQrMh1ypeX5FEl1tSH3z
QAosa6LqNPaCWp95igsbGn354eh1xl0i7i5clwyu5pHVGH5WkgctySs/RrX9cwnt
3mW83zuV3AnbyMPWZE5unhI2gQuNIi1JiTpb4w+9OisRDfucfi/2Zt+kOB0KiHGp
3sfP64fsyZMWeajZ9n8j76wFBHBjIdmyAWwOE/um5ZKIq+PBabbq1mVoA0n2lolb
XDSM+0phi+Zdt3m5LETfzFEcE44e88DM9Ri5fS+SzyvKxQRAHXEzaU7D6Izwe6sL
l9hJfEaOBMzHBXd4waFcy2ppy1J5CR181jbMMFCEhhUsCkzjsfw9gZndk/cFXS4m
r2ermmyJdpovLpLRCV/drV/3iaGkTAqFCUGiEGZ/tOEJg3SE4NtI9lVE596xIFql
q1Ftg7OHW072DVJqLjv/yuikqwyknDmIMt/Are0L4oAVrq9J4NuXwgDRCRgcvtsW
QuVU1j9F8AY3GD7tUQ7GKIrbZpNAGGAiOb/n+z2zFCvTQ38v5oZEo0PJJ7eJUUZa
YFfLSQe3vkvsXPa94Y2PEdkF/6BQH3zWYlrtRBYOLuqFM7ac3P4hgyvkMMEdFY4P
3oaYECatc77Gp069rSn8PinM/QObT63XyepaOZQ6xxJHuOG14xpSLp8tIcIgEUjo
o4u5TuTJI7fqhnkd4YC9ek8jGqcvJQkWfc70QaZBNn+yopBDxJmr4bEl/Vry/Y/V
53foBigcW9mhd8A8OpYgaea+O1vt4WuSJ7WatTjsWpem0tnKStbxNnpOTQ89zbOc
GE6fRTnu3C/NVZWmPPmjp9xU9iS1kRTajp8TjDhCBMwBrBVhd2r2WW1L7EPJ3dHS
pBtvjoqAto+CqJZzpTSbyG1dyf6J4sR/+rPtclLJMqaZ1V8OUuCvwDd1g2S1LUjZ
vWtz4DqPy6UmrH6oVw1uHNQUz+mFmkvNDcQExrSvyPmqUUSEkHAmcDUTab4ve4eg
oKHJ5hQaE0Hu7A3sxaFWo8H9lC6j0KKZNpO/j7N35J0cIxK18iYwSpvPeUeZirKm
LmYZ6PtDJ6/9j/x2yG1R3/ToL/q/6sgW4jTZ4aJohPbWhmpE79tyQ7C4Kn06WXIM
eyz5aEld8c5f2FRZYAvk2Piy72RYIPppyrgFlUsQoJXBSfkQYZ5kAF+Pruj7fqsg
pWoEnINiWXUbrjARiKiPVYkXBscVXc4jij4XTfooz4RODgUKlWBV5UkDeQIxrGw9
7mwF1ujYW6PtN89OCYrBq7nO5vIUREFnojAphHNXG4dUxiiZXYWWbgbebqWq5F+i
yxvE1rMNx/Nb3/KVivTRfYSCD4ck4omq7zRjQZWpXQ/6xOnSU9zwJ8qDsxjz2S6F
kexXeoqr8bagEeJGztSBeRwm54/Smz3o1SZl0mAGWhozDzZ6Xl8B34yVxzsrAzkn
hmz3N3lrqw17nvZ6qlq8+V8LO8yE9ClGt+ctq54S101fE8vXUHCNjBXqNSmnnxeV
PkqjXrZS59ZnbbQARKnzQfv2UYWE++fyEgXcCqxUrRmf6EDxFNRaNv4rruNwb+Gp
jEwujHhiD4bscpXOE+mOxrPpO3rGU9qw1Xtx4QjqSnE4MpZO/ZXpNLYYB0mVUccp
3ZiC+v6D00uRcye2lKx0FDqyVKAejMZW8OYNcElLNx+V6LT8xptFyfnhtGG63tkB
uQdPq0avEt5UeXAcPMoeAZ/KwoxYjZFHkw8j10eABKBZsZr0/wfon1En9aR8CdQ7
Mpj71n78/H978f5hdyNTxiP7YzXlP07mwpLhWsvhPh/rfkaB1Dw8nOnBf9CAYv4j
S7bsckgLWeWUwbA2S7mXYkpJn66apcXU008E2qlzbS/EQZKtp4//SJqP1Ak8IaZZ
yY8Edy+NOGkB/zijEXURW7R25e7udKLBeIi74VRfsmZqIFRR0wTeXWLPP/vr+8QA
feaESGtI8j3sJtq0aWoffuBa2OaBQZwtu2E7Lj1YEd1DqeEpNH49JzAq1DNedXrS
BTJxfR1l8DQV3fUR180NbTFgpwtyxUgbZ3DF0SlNhv+42i6d/T5HHu2v1DdRjEv8
D2r34FxW4D4Hh5eg+CZoTeMqnqHculR8IjpTMwIpmyTe4M5cxiEyzX8md5aS/JNt
WIwZw+YrNmZq5C6sRgKIzjAAqYOub13Ji03VJB/pwQkNomBmVUYK70pBreEF42L8
WU/kVIv/IuZEF1NEYsZAp8k67vT9ZZbsLND6tSS8dIdPqGdlxzQE+CMtu4xyMLrs
zjn3D9IF707bRWZnf3kGPVVKT4JqXP42O3th1mNS2CNMtx7+JYe9R63XHm6hL92+
J+hhqV35b2xwFjI4yJaIogHZfW1C0LfksecslV7d+hsVzujT24En/YV2dimjzhXe
oEl4qg8OnMP8CbpJ5p0Boyq/9OBQI+ZRxtzqWcgcvgD7JuTqtvURgCxMJgvcgq51
Chgy6GImWOMfzhbcpSThjfzoIgUe78GM3W2SiYgk8sFxeGhgOJdgKizdeVhqE1Hr
fn5xw76Jl3EdNJFK+vFfIMA/sNXHqqkqmzfOsuo8M72JpWpSmkPGXNA03dofdyO/
zW3ofX/hAIF/GodZ7mz2TJrtsYPFdAzRwIRCrEen4YN+s/TjcUZYD14TFPT2KS1A
KatJvVxGjY9qiee6Li5DzeXbsulYXHGJJjVjTG2D/ylYV3UIS2u4oPP2wou/Lnox
1PJliGlcW5zfPH6eb1I8Q+RcqETXhskas+ZFDmY7IEZ8UC+hj8/Le6x99xXzeeny
eW9ylP0+Uv0e80mrQTa9a7y0iRWAwJ7nKOYhrOrp+RI1ibq9ujevDvlpQ4ON8fJd
nqkfc3S10Uf72Fr7DXm3PdHoYLdxPr1PNahMTrOyRVGyBTjY0LVG7vbKAEIBbPNX
6at3WoXz+L+515s1gbEVlIXZrcSD0zD+qgTFFSWVw+u6nsWhuUQEh7sV37HCZk7e
bvB1yDASA7Bb8V6OY0DmJH3GIe+2Q1qif5ReK1oWUh7OryIX76obfGMBTmDjKiU/
oW9IlGG/fHJ5Oqg6Nvvbf81l62/z4fi8AG2rV0s2mgfZSKGeEzf0y3qKRpMXgRiH
FdtJU20jn2U61GE3B1pQ4R+naBQgZtU2UenpoZOPZgP3JEYOOMm8tuBvZGWiOunW
fIZtUXbKwAW5dFr4Cp2hV7Q3zvNuhIGPhYdMapsE08nXgL6wuB8d1/S8wGPcYIO+
mky17z7WXCVBjggRqjtFrWO65wDlGHrRxP+gS0RsU0JCqFPNEsnbpgGOSWbLhNmm
LfKJhsJUQaiqBKsMGUcKtD+dFNDAphxGjJHu4c2Eak09pyO2EgraGYg+M631Q4yD
ppZ02qUmHfvo8N9tobJBB0pNjPYvzvMLAY909rcA76IjEtk5tzsg3BIJTUIp5hAi
6U+xh5iAt3KCedXS4M20x7dZe53iV/TuR1zCkDkS+xojrigp2sKbY4EZZZznDq6b
aLuHbzYfdxyxQpqe87k5JHPpClxNz/K+vG9xFQJakoo9G+iVO+KypMgsaGobv9fg
vedj3y/9vJKEsrq0LzBaItVfur3fhI4Eu0BcKqm2dKzz3vW59nx26L+xvOWUBCXt
L2Ro0AeZ3FKmAgbc3H2zwkvvYP3SJnjmTJFO5EkMHxh3/cSG5/LiLI1NK3ZpxgXX
1jGNvepmbc1DinmkDtgClZZUBqqoi0C+pEMVuHxe0FFx4vvl9uVISuMZB0RjXDCc
aXy3tfhA4r4c83lKuqAL3q7THoS984bVvo77zEzsW8A1NMFEIIqVBvksGv7BFuTy
zfTlRoQk74bQHSaAJhahPp4WqAg8Wn6j5LmTSQX9tlkA18gKnxdKZ1lb3wJu7NyJ
JegJAi6mbK1Y+jH6UlhrHgsabeycs14Y4uDyH+/svwhvE2l2DVc0OJaPDhOTRhTJ
KXAuHdx62fcn618JzSOgY3rnkPZ+Uqmb5Kfo/02a4PBJA8AlJkwr+Tz323miDG9x
wodzZWXCNU6swwHmNAiQ9guVU06P4X3gxFMxSJqm9r+ZOUknP3bALcWBT7zvDIvd
ZkbmFwI2ra6gOxxEo8TAi2B4xvNC5gD27W7Fm/JuNjmwOr+B7dC33S37LoNg7LmA
TXJ+Fa7d5bbkFCzRW+NtyQyZLSGnmsqKs/hykiWM2FWANn0GFCqbMgDs/0UtGKnX
sSi12kT96HVYAvMi2yJFhWg/zyHZ0YQKRfcc1hRPhqBlkFVvGWe4yoSVKtX+dZZ8
og+OHaVdLItf0J9Arb2ahMTaO24TPIHIVi96slmoXCsrVebPJcoIdYuoXrFG9EOT
Sr5N71LOxhJVXWVNHtiYnEjj6uGTwm5FpZ33puTOU2a3iEwAcxckeOw+9GGkvEZ4
NY3OXeKRtqc5s3Id1guJx/Mlq2N3nrhjgQTvnBx5oOgpuG9M0auObtkh93I5C5D5
tadjY3qV20StDuCJnCC0J6D7qgMNtzR71M9GDjPpBuQSWwmOASDaucoHFrvMMnQq
U3gCZKwVYLtR4++Do7fmf8hRvIXVgZqZ44eltogb687w2k6Acmv+CMUPUuT0yypB
IGe2Qn4ZxgjhmGVb00Oysu45SJ/cvjjRHhJNK+U4wKTN2PJMyeFhqVG4j4KvnIhl
5EqDGypSOs+9d51KxkVeIg4Sa+/smsRZSJEqLU91+h9jO6QpoWQO+qb3bZ4hV71i
1uJnAta8MXgVGaeIchFi27ALGBeSIHmqA4yJgDsGE4k7KnKAG6tI7u5QB2nVzV6s
VmdzCdDK5xX69t8D5+Uqt4brtdA7Y/S8qPxxer465anYqkBIgmT5POrFAsjHLbGa
+KbTDV5hvnHDy5W2JxnQXJvSakCOF+PRwpGtgogBDBzm7ld8WrfH2qm5HT3clTOa
J1hXT0f/1uH1uTDWCx1QS8BIndphakIifnbSFc7sKC0utH7ILl1vRv4qdvOpBPwl
gzPTp1n3nD6NIp4HfgLpG1Wio5E4Q7DdVWwQu3sec8/hmmAvZZz6smwB+fuBm0WB
4iKS4JzfTVH91tqqUKSAc7ZxnO8rrF5SK93xx8ywsRJMIX0iiUfxGLzgfNoGeEFw
dNBbeiomE68B+3+3NuadAxKuJ+7mLoIIIQ6YjdqMJeP5wXCwjru38RtmNPE+JbVd
3My4jFqWDRejY9KM4XNh7fGrQhvmsOwyepoHs7zcl5lQ7hJ6NkZrcLYX9u+auz20
MhSZSuaWfMTBMreGv5cpnANmAsnAIjFnY/o6ra4pHBR4QxlpE+Lb8FdfpgARM/Zg
fjsNLQbGooU2dpByGHbfcuWc1aQybrdmLFRkPxCbgSUj1umG/x8EDb+ruubpGqK9
eul0puHVZkfKgpOVkcyp2n+de8/Uu/X+dk2tekZKA9nWs+EOVMBTSyFfj3Kd6caw
rFNdiO50vSOQEP0ZNm0RL+YMu+oSiXidZ4uwzeZpJSGDKB0YNCuTN0AvSHc9Jup1
Iqo7SDO8cvA7Zak8scGNIGKSm1TeSGU+lCn8DeBWt7nuxzZttAaMwAmQOweRxcrG
LOqusDmuWsas6o2XGTidSz2BjFRiTBAuLrPSqp4X8OM8++iFCdUC5elP2YUnhXj8
tXPZYbT7zbsA1x9j7ub7SMvHYUv1V06/LWEvlNuLG6cSFCIaXAr1MCHdZNGW5qAC
SgilfdYy5q4KPtBKCHWrjLtn2x+AfWl76urMnZvVjKdY2FOEjB5xm/jAUp9+Bw6a
RkfRSSEf7Tot4mhUqFX8SgWaPYUHJYui82o/xAd0J2NzSidtdQO3EBYrF70LwmXA
IuKYXpVtw79y4XRoxrKdcixhCwcR3Uh7Ul3ZhZkJ6au7TKTm5hH1wSDouBFd1HiY
mf/4bdcj1985dlLR6AiE59c+RWJX4Jvv0ekeKmCZJOgWxauyw0zMTvAp5OxLCeG2
3wQs3apLXWZ5PI516ewFH/p6oq1ge8jatpsYjRaA4sFqxeZ/MjNdi/mewVZIgrR+
cDLTxjDPHLCCf45kZibUPoD2umZokX7pg/BCduMIRtcD/xT8b091BxPlHLasPzQh
evH2mLwKprsJsY6qyrNRcbgLNo3c4WO4PzTyZDPnMDX+qjgpC2vuor7vbfr5WJ3R
xKAhO6xCoprzVbUOUwQYTN478xA9/ozlYLmZdDQozKAGJevR5Sr7vh8HaFBMAQJ/
n+4vZmi+0criT/4s+HYAbzY06gAMmA4yUMN2Z7ulKVYkEpDeB7J76fPexqwjr9/h
cNd9igMgqCoN2wTc+aDZvJV+px9xR4VWQsLppXgEb/T1FywLSon5kGBu2JLkUG+G
kRlzdTG+m6cBysU6KU//RaZe5tHmBDCT7KsTvc8jp5HWYXblIT5aDRs3NomFCuvT
08NKudfbHthN8B0Ds88tGvKMbGjc0ITLKtkFTS48icdW+YUc3/1GK9ZMjkh1FlJh
lze1Hd2ShM2VG23i1TMIO7b1Gpt/I9UuCXRYdm2eaCJs+qIeD5RjMoLO6/TWyj+w
UTbmW9m5oHzVuQ1hEwxE6RFmtlD/JT7QFt7rfCzMupRhLFpZ5VhA61aa6NTqB59I
8D3+3/Inbjk4sclhJD/61obIqJF7AXh7hUtnvVzNfRHVkCWuYyGWT/UY0EZrtsaU
Iow9ntYCAGZHPmo3g4DEFTDHF4iqm6kLE6qHhfjygLK1/rVZ6mmuo/KGOLorBNLr
QP7iOVwIoE50gzc4ZFCm7AC50K3P9lwWRAB3HtzoJ3mvSyXY3ccNcwryRMPKQ4da
7d7RYfoZj5L9/YSF5WxMftuSXm+AineU+C4BAomePqKC/fDhjC/gacYjXOJnrBS7
BoG69MwcucAfNT87MhdhsJFejSaEqi6OptJ54kVQXoLCNEo7zw5b2X4B4Y9zzZI7
hihgWcS8WJVDQmgkV8JgUYKqY/BkQiZBxDAbr30dMBx502miS2WW8wZmOHXyVcdX
qw5PXsQ8HWYVHMtfcYYlvjuXqHNhQ7s0lNElfR10EJjfWc9RbjAfHtle1vNk24ye
IEIRtVT13S5Ri5ULXRw+hz1HInBpimGa8doZr6mlzAjac8Ov+VbHLmweZBJskLgk
8rqc5vmMjiO+1NpDePSj/yqbcNBUEIJwNws040+ihAQzJeqzCOJdQgeKJb5O0JUz
378nMk/3OsSgpUt7cavu+7QBbhWiwzoQNaVpZ9lYV8x9Alp3iWVqlvelsZskCf1C
xo/WcJHaYwK9znnayhDpUglcKtoSOq79au3Xv1ChDUlBgIU9pB8EnYnGlammbB7b
vGG0uyc6jWvtB9cXbwJHmUmARjSVKl9j8TExf7ewgkirAx7tZhsLsU11/9XTtSTO
BazhDgr4IgVjhC8Y4jXKd2/MA4Uq2wX5aHnW1I2geB3Gk1qGePESiWPdmZt83fa/
F5ih6WYoSUveun22PQLHI0YxSSfsafwhvAng+yRcuQ1l3VTuYdz/Z6mR7adsRbLK
IGt39yGimZ+zpw3ktUEKPY4/hIEqRNHIAnHzk0G4M+SBtUJCNVLdOBS/84xjm6pl
Ak27dGI3gZlS4MqR69HzIczuVSmzQugg0MiZD6WsTGvbSMRjNK8ysHQBGQG9kVM/
Pu+paMxsdjwy1e4rpryyusnGc+mvMaoXyRMEMyDJnqAIDw4wdxQskQKOLDdVRzik
NFDK5iOk+Op5MnzPPF11FusyxrfTvaA+nE1jNrtXaoMxPUjdCTfjV0/bNCKn7/CI
bpWLxCHCV5uXkndlohL/YFW1k3GMUC1jHtmG92E943OZS/L+ql/pbTkpd0EjoACx
Jj1sJD03CwAJR6XARNs4lVkS4uWplJIP3Hd9E5EP/wnBsvCMdPsh9INjlBh2O7P/
QoSEdTnYdLPjgClnx4b0CbaWXfXPZoWFu1ze8JP8r5dhQ363NVHRu3kPsCx+Uvu5
/kHlJAiZNkKBP2YRCrHc3VVJMIKKhXyxPFi9I/9heeDOmj7CCNpAbEHuTEIJgf4e
ReQnPP/gcS8B5Fx+ThyByFTXzMLU6q4u1flgz1bmNHlh1jqGeL7uW9zHBcZRmBNC
H1/xDyvmo8PsrBLZHmosYSI00DS3XwyKS3MrMAB9J1p08IuUjmjWLlLPhy2jsO7o
MgzFMhXtZoFuvEnOVSdIcE/prSqIqGrjmJ4hVR6tpyjHEdtwrzloqGFAjlNzgBq+
d5RHOeHQnHlASpo1LTJGIeh1Ku2yoLGW9CHRsyOXh5nOpgFfrrVjlPHmsI2bT0Br
X9QBspvMFqRpyI8dvRacdAXIvKhWufrTjoDQWlyp/uiMRPLt2b2P4bJV7fbjHLZE
j8NPvzrnfgARjVxakzp6BstRwyFo3p5PPzOxlhgtfb922GqB8zDqkApfPcugaRuY
TrmMJfSy35cQlTY8XEWnj3aT1kYfwCQNFuc2hs7KkAoiShI4o/23AlXUG38Vw7ab
icMDtH7bAqrFp4jL4HFRHj+apB7B08hU2Mfj22hmFVpiDQIBZiAQxo4DGKkLQCIj
2ShPWu3yS1nAPMBlt+GIqQEqPliCXEQTyfbWPHh7Zypc00V6zcJR54m667Gz1+Wl
PUceFXwPS6VXhVupta7mUcUOkfuUIb9cyJ2DPXKhLkVAyqWOQeZTcO7TA60YFKmb
sI08cre/X0A4WHYtQRJTQG471guANwF5oBMkwnCDLlAwCt6cOnDu/qdPhkU3u+mD
fnr8V6JZEhmk54EHWkJaylXMaoujjRq4Km795P5OAsLQpapSRsdKlBBVcjiAiCNC
8TlTYj78UcXhZuRtk/VhX6Dr4tc75Lifk4Oxl12vIp8lxoAAP9r0nf3tF2eANXoP
LqymfwdJG5UqEBiEJFbI3B+dZBUVXieJs5rdJlMEqdgBVt6sw4CMSWFlpH7B2CZ+
JWskVHhOahTrsDa7EotPpACkahYYB6y5fP7a0ohrTuhq5s9Su7xZWOCFgk5shPWD
boDpWPCzGtrbtyo7jlgTP5INUzL+rIXMPK7d2u7arUv7qMfin6/srWwQJuBIqYb3
lvg07EgEmL/6UurmW+Rnm3lyZ8tvBNyAY/FuIAPRTaU9qxNYwF9Aver3sUzMz2pg
eLpFCRmBtOHwhtDssRtcgZB50e4swR1SNo47di4NBaiuNf1E4wTkbnVks3gHxI8q
kWLq+xoWpTW+m8Czb0CfhHqDpoY11Eb2GuEB+sW8HN7VCMcP01Gjb2SgidgklU3S
3n95kcTnmkuhLHNJrgeqUgCYgKCw/bMUBVVo7Vi5r5aphqZQ0SEFJ0Pi0o0k2wKr
U372KIerW5l5KWNxx61cKOK7XeNw+98o49vNGyEv+AFbC5fPlI2C5tquA8hnrjVk
+JE6FzMILHtrfENzzaRkNECUVy7REdo2glTzxnFWFkPTRaYUZ6OsXe7YNfsdNtMP
hz2ofPnLxe0hPgjP4J0lxB9eqBDSRODtF/BTRqmhn6Yw00KV8Yrhok4uBaZ7V6LR
mgGuZjseZuE/bcTAs6Uc7MZ3kU17B9gPuKAnL1FyNkpXJ9MJNn7rFR3Fphu0agjz
XyjiMpKSATXwnsXrafCn2etMmU5PJHCHmbIZnoubx/U6ofMkv4ZNfGmR/KKy1WEz
7TSSZLfEkrsLk0pFlPFksnKf5j/kGCe778AlCbU+ryArwGFPFwReA2XhUyuIrGQD
9MHvPOJ/LK8WZgg3aUvrOTPl4EEYev9OTCTyZgMIML+jIpB24yW5ndtIOSlkQYFc
OGMCvaVUJZGe/NmPWOBO6mUw8MMWBANKrJbWydMU0bAj08faCw0CU+HS2PYX80U1
JsUscGfMvGsy+GXwnfpPONiOXlpBL1ImRs03PyYPi3ew2xD3rWBf85LgayXDgPmT
7+5XdTvNut8rlrwiSRa2EAjnQVDgdrtIsKne4Abz3wwy6cWMhLIrMbHgiDaJXzG/
uNUxHtHEvwxn9NI6CLiu9u3vUnl6kS0aIfJ992HcSKNNJRf18KP4yBPR+D7Nb98g
5VqH7zrFQ/vXGc9sbelM2b2WutPV1E4N4OaLV1HehTHZLcEzkpQ/2ckoZzqtdMhh
wWybL8ImFx2/m0anBM9HlvYaW5fx6HkVO/hJwK8W/dnymMPWuWuhFKOCrTnoGxhh
ebo+oE7M2SRkQsjS3+VYXiq7ICU7Jff6bXKglocKkIzK7FEmWK38Lxzhm35MzLpo
rqYpo//0ZWpZ6Bzww5e5ZaWFAXabNvusJf4JD1uxNi4Fm1evb8qP89fcUugv9aL2
J0/NbPX5sBwoMBwWt+/c5hNGZzWf2Mz3/z989VHeon6niVQjZSfVWUd8nMHQ40U9
nsHl5xsVRvhr4UfIyh37S9wv+Y/G4BTPiw58Vr2+zZ2nbg5jvWFY4vaPKylFjWX8
r8x69BRD3TGWK1vxmbTM6uAxWzsnvypIbe16w741OgvmECdcngEo/4gqYTh3EZGo
9BpOPbZxH7NkicSPjGSPHGbLki++IQsZ1S0mn2Qudev7JE81kEbKQ5gA+HQO9dQJ
qHhz7YjMwsm0FdSTuzoqKtuM/dqwDXnUxVLqBOq9UWFM59zSH8F0CwHThsGlhg9I
n4OX/eQRnnLRhU74GfHw9d5U+Pvi8iQBucPm4bXWNfn6paNoNw2M/UJIcITgERDy
8+4+jpHkiVYXlaVwQB9fpB1aAYWPuujfKRpWQtLw0SfMy8YVEM3ROyrlZvGHSt9B
meiXTYspmknr5IUyYTRxgXpdO5+DYjCn6MDsngp9W4xFKzLyhU6WLRiy8zXDL2IW
UtHVblgkAKoi+oNh+XbITTUVv6U2SkY2R7ISOlylNWEpRqsbF3OSIGj5kOLoSBIl
xRQTdNiELA+LlEtTRdnEDfM/uy79UP88+4Ca1kTw0CvlFb2YnWRkhmQ54ay2EpSS
+srUgP/tGn06kNoMM333l3k3FcnFb7E6Oca6VVqmBMb0ow5f3KZN5X7ba88aL4A6
ulAPrAZpp3IgNeBMyESOSfqeHQ8hyoExpDUgwO+xd4wQJxYLu0QQmGrCHqNFaRy/
4RuM/foPJdtx7lWzimmAgATL2VSxirN1diBj31fdf21k6rkRHGdqPOS4aJaFcRl9
iZyhxgC9X5+6A+urAoS2ZS+ySddTBuyCwgn/cYGV3bUkAeEvZY2sPWGGwGyeAbAW
96awe9e/4G0Ec0zTYasjSpxefEyK40HGhPPIYKhRKzjGipBhuYiTMXj+jPro2a4c
NAXw2roaDME4+dnUPhXiR7i5Znj8pa1KqoWprTCukQYFjRc9WQwjCsaBdYxoVxKb
H+b+xcbis9Q5/OiyESq/jdJSk5hrNaWPh7au2PgRvNj6oK4Y9/FpSE2p27C/6+I3
jhWjJZbea+M/EP2Iq3SsQo6HA8Kg43umJhz/fTC42IuPxLstPG5fUv7Xw0S+7ku0
6u9ztxioKVGaqJN3eo9lmIz55m78VNbfxQGqU1LI9Q/iPJdlsl6ALM2WA41B5tOS
86P1clBn+adjYJN4ekfHHsHYA9nSvL5klHoNBT7VCYjEC7RPqb4dkY69Nk0UW8I1
3xU+4QPYuZvEIYSmsTzioDcCcc05fk7r469jb9fn/DBXWU6IBvZZqVnqqtRLKuWP
8oM4iv/FQUcwq+A5q/q1gMKYOyudqPaoGnePn9aacYzRJx8pU03tDSqsOwd7Ao9a
MF5HIP47Fl9b4ANGThUQoR8uWaynhCOHmo3zSHdaSKZHEXg9skcXiBa2qgmd6kB9
YfMMGC0S3l8JAWZTiVISh9zfOIMKDRSnWY/f7N/cgnYaxUIIbKy4lvH/eKZEpJMW
WuyKaOPA8W35wxnmdZrOpW+h3FY1rjq8uLENCQkPiN9xyofKoEIiCub4+r554UzM
juw5ewhs0TungLfN+J44QtJnxPEMU0eGCJW59VkmLSAJwOXyREMpG+KxCFHwvCeC
1VDGkeW9l5NGlucBCttkblCtDsTvq2c+Td9w33IoJlsgef67KbLasuqZQnoFxffn
yQ8yTI/ykvuE/+g+6UpwxtIBQT0rcoVuELs83OdBInvU564XSRpIECNFseSKRPt9
MG0ZvR7QRRto6/0/awIfw8/nSi8NIOkDolx/on+tN30YX+OTJdlnCz31FJzDCJQr
z/vWQ9KVSx4xYRkhE/q3zaYdSq+D6JBTXbj2GgMaXKml8aXT5/sKGcE+qSlYdacw
1O0rbdtvNt17H06//f+ov4IOE2I76FcPAGGtxC9pwdrnQhXfNKatbLROmwEEuoz+
+7jihwm767BkkBP1dtakFAFxA9OkZ5thDjwo2MA2LYvgpWawCPKMMCOs1RI9Nq5+
gNSbH/W21bznONPpz+nXeCkGi2ptqm/DoRN71NeSDR+lkpM96ehNN35t/i3hNJ9s
a4IFM/6SFhtJevucsaGFqKv4NV3CmPxxUGMLtWHVjpiqnqXXYj0AypqYgihp6+Uv
DrH6emKXDAX+CbwQAfOz1xE+L5TBSE80nbiilrSIhQrDO/wWpXJtNTULJUlJv5k9
P/mWS2Nz+FUirN+zxm13MRFCO2iwqHOtFB6UgtJ7E39Pe0s1+0UpxY0tvMraBews
Zr/xeiGjJP5mGswfPqmlVkhuhEPaBPKf+4IBymbWu3RN3++HwYMugvsoDK7doVZK
R7MSARzt9PUxMO+hv5juRbGrvouQf/+cObPFh1pcsBwJQ0qdO2xDNbfLKRzXlNSZ
0HrXhAm9ECzhfL+MoKelS8iUed8EdPJsjQ/Ywoi32R6WniExT97PwS1SM0GTQpgu
5xeEz6v+hl7Jt1NDnK5GJgvtT9/gyZcHH3Sgmm7jETVl0ZBRYrZ3tEt4hPXbfjjt
g3yoIcmGcjXS21FBS956aSXe8svhCgV5OPsS54xrh96wVALemrrCaBBdWF/t/u4q
6nEfhi+QtblyAmgV+2hKwITeJFhjoPsJX35R5wV3SqfE9EyYOvikmZyhAvoQPfBq
WHhfw4NdJkiq/ZPCCJ1Crs00NhqJJB7NS39/xQ7HXsKrpn5IUBDXfdHZeLucePEm
ggbjE/RO+G9L0YVO8x+Soz+8fqfpQAVkXg6sjYigbFhLns8CPwDMYije4J992S6P
/zgSXhQ/k7S7ZTkcbKX1oARPg4zF7jb+EMQwhFYYJN0THzifHOol4BkaL5gGkH20
pSthyGS77AyNf3CAvWY7IbjuXiVpvOes8ES2/yq0OJ9YqQx5WiBzOSaCWz94ZAFn
jjpXa/dbLBvIDv6lOEttzAPFEBfXmUOorM/Duuxm03VY5PK+SwpwmHoP/NHOjY6x
hHZUqMA+1VWqKbFcO3iDJwPX6+yDxmCeg6zXPnG2FXEodRBaDZwux3UqX0B1pSNc
bKgUJScDy9kCGAzzyogtGZ51Fx+ZZw+V8ovX3HSd3eGAfXNTwk/HRKvsuSf0rYn2
WnN8pbS7bOXOvhaucl2xLmyKrCBeETblpy1XGzb3PoLAnK2IxU6aIyZbscbP1Nh7
zuU5HgImEA79DWFJ+FKB/RL4dJ108ZxU9185tw6LKEI441b9lxI9+YbXz+o1DjS3
qrS+mOhG9xvlQeK1LmpmlzjduKjFWYvGZYGkTiaAF23E6vV7ll5iNzD0Rp7nVF+i
nb0H5qA/TX840I4+Mq4gkWAj4xa0hB9uPY5LKDInrCK2YVxXuAthxuUpKw4YSit9
lDDK3w4BjnrhBR8NZIE7/G6zv+cmcvlipjIyJZAEkWm5yX/uDuOVnBikc9j6hr4J
M2cS2sas0FUUQ/+jxDJgN56ZW/+UywORL9V2bsNmd9KreSImlMInz6WrnE0jB6h1
i18EsGYjxvdYMmEqBAlUlhndJ86TGMofRhrb5oA0WYh+nBSEEJM1w0UaDRV8GukC
UPvKstIAnMY7dvqKZ3WU1F9ug3ox25z+eSueVq7zeRl3yMHNNqenue3qKHAuoDRK
2LerQmWyuOQz2oqfhhWXlb8lrS5X9z5t8UPG8O4GHkoCnOpzUN1MA4q7IV50jJvA
qJZzBkKF3CskhHLfnQwSFEv7E+9mom093XP6C02Ew2GTog0GChjBa35sX2mbubjD
pOtSEkDmwTensUR3hxtVDerd1ZuToE5jaRk6Cc44Nrc6qx1eBFighyUCBeMnQ15f
d2vi3p/QBet6EFzXKuBWn0Pi5mvbEJXuwYoSdJPBdyVnpoRutv5RnvqZehjAh7CV
30eWAc+axq/koDDa5eALMeANdSXLHxiUCAZvqEflfgNi9kmufbZph27jBwUvakv2
Td8cW3mDVfHVY5oWsCVfi5sMhIk6OVuOIJKefm6L//PB/QqFIgzFyhcJ76qf9RgP
C/sSWV0N+EUDsu22mV9ypFrjoh1GeEMGQ2Y1vF8nH2hE4t28QmRnDahyjjBngSs0
aesGvIodMrdZ1aZaansINUhF/bEAJcRlNJ1PJRhhUKUc8WI1r/HmX/ZG0feBpe+p
d1PYv6NC1TAIeVne18V31OKHdbTnofAzZy9qmGrH5QLB98qf0BXB0hJwEzdrAQhQ
ZfOuxEvQ0ZQ19D9bXiHewx6VhXYm3Q0/juYfHj6HiG/0BWw6xL/StF7EKsFpMWkD
4q++aZfeQL2cM2v9k00APC+Mv05oOmkVnHrmUAkbnQl0GofaM9590OFI0q0GK4Tw
awx5/6EyaE/uEpgJs8u+W08dxepHqYBGKDz7JzDbDxnXJu9d0w8/wuYkz+m07/28
sSiRyilZzEnLtUdZH1iRELLRyJi2S0EEPLsHyEzPL+sZipv8v8DrtBO6OfNxW4Er
jm5gSkvQlPZaY8bjNeu0hQ==
`pragma protect end_protected

`endif // `ifndef _VF_AXI_OPT_FC_SV_


