//----------------------------------------------------------------------
/**
 * @file vsl_sb_report.sv
 * @brief Defines VSL Scoreboard entry report class.
 *
 * This file contains the following VSL Scoreboard related classes.
 * - VSL Scoreboard entry report class
 */
/*
 * Copyright (C) 2007-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_SB_REPORT_SV_
`define _VSL_SB_REPORT_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
iAQ/YERNCaG2JtVsWZjGZtkLPef5VQwfo7ftzBJBCkueJT+Fc0jsR0++S02SngI3
3OqYf4H/dM7rse6rYigvg1xPYiYVgyQLuVddkjv+3Ox5kKkrNA+g8By2RptNuGF9
nn0QKcKW7OUL22s2TrnIw5mJ6h4kavS07GD45gZy+/aHT2poYZg3am8PxyQEuWlR
/7H6kk59zVTErtZkuVuZFQ6vX3/JesncaD7/5hn2Sfg3inhLd35l+3zLGX0/zgbS
iboH3ou1SWpAg/uLt/HFj3i5Vo3NymYOr9dfwbOhCcT7BsSODpb98zbZSHIk2F2I
ijgh4whJXvCEdQDwISIY8g==
`pragma protect data_block
1+8HM3m1o6o3seNg6HimfLx0NZYAgscy+g4oWnPOBdSAO4ZmHHSgHyiMyzqpP3Y1
y8egxRPiMaL5GthIpw27OE1RD5i7WrvYQP4Uu74pTvQr1bggPo7nonoGWXKu3NYQ
3Dq9/xY/Ypz5yQog+UzSs6zo4vk9HNlKR3Y3pT8eTDS4l2k/nh6jyLOeibxV9vIw
pIsr5NReuPvqVdpJfEFNNrAMV7PQ3wBgNjv/iRAOPopDbqotLErAHJcbK2VaWkXm
bR4jsMU8wNJ+n6rfMXyz2iP1FZQTvHzl22sZTod9Wfmkj9keZa/YXfx/FG0wsYnC
VbXtTmbxqfkeV7tYLJ498CgzKwhFkslI4e/WJAp5wlJrB6pEb4N51xADKYIAChWI
aw2FfwGBsWBGAHMrc20xyBpX+9IZU7u1BEBm/SeZ6MfWel/7xZKiTrnMz5Vkmbb0
txXo7VLymtxVKIvDlRTrnd6+Fdcmg0ZbVCQQtuoRYTyxH59RDTD5hWzk7CQuupSk
WE5/SWOcMt+eo9VbH9czLBzdMlp/ztInYDuOVRUWqF7UdxQ6wpXgd2VGqFT8SFi2
4LiV4704908efP3AA3VYSO5QIt1+xGK01E9sK2TLf9F8YlUmxxmdKrXhr1sP3cIL
DFpDtcjMge9tYPk5hTTFoXOV9W7GQn8YE5yw+cWtzGFuj2xGJVI5+4OtAjvwfjp/
b1XuM2mGLro0rpkqHDh53azNZkAo3Pd/kVJwcqucx8Buy3tfvX6SQJaoiXLg3MKd
DWpz/VsT0Q5X0peWIM2szDs+RNul43jX4ibdTiA/KKLCG8gV7n7XwWIoUwtTb5Ob
AwjCcqFG1cJ7v9aJrvggkJpZtgbrj3cj4w4uzq3vrZaL1r08m/odxaG8Nty9tX8O
VRTKok84GPHaMPddBd1OmBggxGPSXxkV3hwaH6v5akK6C+fgvTaTQnnhUvHo4hPX
fiVfrbimbOxYrDdE/NUcRrIk7iSspRsSYd/MEWabMUQC3KJxkRVdmPxD49+yTOwe
XvG5sGx/tDBFcWCBmC5IxWXwPybBYrm++67TF1gJ5f9hs1+ZbPpTUYpiU5eca+0h
O9JZrM54rWoowhinmnyUE/EUHS3f+171IEe3UaB/55RH6jOvhJYVnSh7Uk6gE+N7
N5Tx0jnd2Aa29OKFfKk3Ur1aZTeZ94u0J15bAENKoQtpmlhRWxeLmWdMsaxjv0FB
+3OjYkilmThfUWSpgg+9D2I4NygDnIhvsOSPmoILYy5aNjN/rgQXvXUV2/mpKKFw
KPzGTvyjtTILng816I5Nh0Yly2/FAOjaf7gxbhO06DDeT+9SKyeDw3iDwoaJujte
nWUjIkJiv4Zkb0k1tJBD6hGLaO4nRRqbgXdPHyTEzzoABhsHljhSbPWbPnoo5/jZ
PO7KYsbRDa6S11znyx03vMbKjp8WZ0yn/ZVth0cvBFTO+NHWhWjrpIz0nzbsmBZE
ns5f9pHCPRhh+SRR+hYkI9oECis2asCqtQ/09uzlhFHFCd4k2rroAz54oezcA7MB
9054dcIn0Xl1AiW4uFg0udMOHtHzb4D/cJTTE9ceL80m+fXvuQhU/5xbmnU7HMi8
xWD25yaA/RJ+alF88gbrIbgQvL27APyodLXHUuxzj8qYmxJVGg84trIJ7hEnBG3i
7iuv2FeXjHfxP5ToH5qEDdzDGsOJpmavw+CzoSf05qcQEahi10ORGvLGES/ItzpE
DbGmtrDzfmgDLeS4gK0HzhPtWYWQbxWEZDLu8zrOISUUumOLfwJ6cqROK9SbB4mq
bxTsNhQGxtRLwA4Ok/qwLmBuCwrCx5V0iM6vGw2j3E1FyLEW1ZYT2RLR21z3Joz7
PkdzI7R2+nXxLve+4es/OdR9Hd6ixZDNFDpX0Oa6jMayqE7odp4hz//aR2IrS9Of
67HeNgvIXP5KSFQ7DRTkxctff13uOwPnTAZ2pnPmWlFrW7s5DlE+ClVYq1uPlwLP
XkhlFR8iBsypMEQHScO2uF/tjtJgrtP9P5CPsaXhMK6U/oSTivD1vXijUmp9Mmmx
D9yukBELbsS3PyS7u+lOO+cxWuNqBYsTmu008B0ul611AChSgh+z3kdtCY9wMsyE
c+qhLM8fyaIn5rmQ+Cp8dWfr6m9M5Y9fTEHbmM/4ZSJmtClv95BEcXXW+4UzehGr
GkRzG8Q71BG41eZACrgDVIahl7MRM12TZvjKmrD1lDZZFxdztSsyJxLjh0+6mL0X
xPgD4B6zaqRiRzSChvsFkJLTchTTwpg7FilM/ZVvH0XHjlkKpUzkG5xabvGYZIAi
9A4NRLOdEsV6XK/hbj6T+pfUrAS/hVdi+lHE7aGhf4O1mU42m8iCCYWwuXYhr730
ImOlNJAorHeLLnbibeOXPF3wubjsIf7160a8JB7NxwjAKchVI/l77fk8WIe7DuXc
C9naoETDb6BkeM7mguKxMlHwSczL9MdIhpftaKCe7udN81PhuCmr3gJMNReJL9UL
XLzvTQ4pFNRSSu6v9YCD9pghgiCAxZxOI5bkm0b/wrL1+s9B7TLDLJKW61WZNDMT
zo2kp8YsbpqSnabnNCZRKO9PKAUbZn5b+R2X0JJ7yKohCgvP2Pcuqjy5SdoUZ/u+
wfLvksv+WUqIFvu6cgWgLF6vbbB6jlo53t1UBBcabEgqaQanP5GHtNVuuRd/SVIr
G/zyBJYtJvtJ0WlIkpci3KEKe9G2tBxhbxR8Ilrn4D76go0K2IXGetVjZQyjke+7
HfeZH9gxThw9LKz22Y2SO/usJicy4yQLdAaTRk2u0hCYaHqpq+aVPIidohgkb798
uoYosLb6ziObFGH5tXoj8RrwrJafGtqT/VD3SPIZLHAtWK+ghrABFYNfMRH4pwre
KI2QIaEkEMCtjFijjo5pl8RfbC49cQzQZAd5COTM0VcIDbjBaFAZRAVOBXbEJP0Y
XZ7agMZznjpFHtsbS0aO9s76RuHXBGPPplt7wscyf0yvLfGSU4unG5iROy+gPB/9
lydALDxwgOP+u5vNrwAThM//SxKAHp2ZcZiH8rU9T3kBicj3zhzRnHKiG8f3FkRj
KVq2anLwuP3LS24GVdr629Tc1cGSq4Xe9d6FU+yH0PAE2FSy9LnWZC7aaB1pL/MJ
UBR3ddRuwHo2e0icP/5MkOxYuZzg+s5r/BBs8IwZDc2Rnl0Y92q/PLF5luueiIe0
KOes9mU49/cVH26EGU71aRJ52vBWQawJQ3T/dEQEK0jMVrDLldVTH99GP2rIwJwa
kP8rNKOtZLVA/S0C9mje0q5UuheeGQHSeGEeN+2cFkcQSDoQFmaGBx8ktom4/Xtq
Mnzeyjnnp1G3j8MbgXNK0GLL4s9mhkUgDmhOQQDT1hM6GIQhcnGG1xZpelIYOjf7
d3XqkCd4psBKYMHkupgrkAkc4Fn5bUUCIFBa1LJMHYZuiWoj6vmKMBB9XHL2VVLE
3LGKb0mkDEzySNDLicx/qMVjV9VFZyQhx7E1cQFqAoA6HAWlZa85NMSpLg3nKn5e
TygXcfHQ8kGFzwIgZYelmWFoOt92xpQEzucug46hS7oqQvzd9A7b4etWJwvhUXtG
2r9gSwXDHhkzsFuk9CGJpW5DZ5fgTTao3lsuXaiWRySo4z3JLKIe6qeAyHa1iall
EHEHmcvfp65eavhw+43X/5bJE2k2QbjmwhZMlNnDrmXfdKQ5i79V9oOzDDvwtffU
m/ZUGOX88LMWNFbipyinsQry7airtIVGltZaAtM+HX2E2/gERxED8VUIf/2btKIo
Z1IIBdaXqPps3Jon0bLxD11qL3bjFICb9G6+DiPrta1he8idj9gaWgZ7h0Nvn8qp
yJmwtDkCxBMrzmdYYsMqz+nsZ74uBQ6D3OfgXymUH1o7sFHWEdRdrULnrrzE27YE
oyWQgSj8oPoqN6+WD88YXZN/kyLzGJ2BCSF0gFysfUaQ3b8HJjM+VpbgM4akBRey
efBTO6+iLS5LKIxMcvMQTaOvG9ikB8DNAs9TO5tOqoIfuzYWW3UtUGd9VbhuIYUO
AltBKMpROSB5cXKc6uyK6A8sRnV1D6ITRJR32nPzlXjA4XCLMgOXYKR/+MVmYrgU
xWLg/3eN+Aje+fZv6umd6A70SMiIC4PxmWZa3kcqIRi6HgJprWC59UM+IvuI8PgO
JZg1Xf9X/a+sabvrhvfoqr47bglwj0ytOgsr7zpUt2YvEyFiCpQ5SbXMjIvT3mrV
mZfsoC8nZFiUMluj82bdBol5Taw6K1jCJdVwLBEchXqJl3+DtNpOnT0lKP+h3/qT
6QF6+UY3KthQpohhQc+9+OuiyzfA1gh2Z+3CiRhoRsacuA9Q3YM+66gn5MvZdIhl
N2hoAV48DGXhC0OlAwY+IeE0G6p5v9NiqmpjxCaCCwwZOCzezsN/Mky6EtAMivPn
eLVOHJPY2LVH6HfEEgtDBj2/NrbFmR1AQLEZv7kZT+k6YbQqMUTCMrrAvIWJiAnl
0wUdGt2W2rutAQ0OeDJLbSbQItyf8xeWi0fmfbnPEdnBuJBIswgZAqbcL88+Bjd9
q5hiloBbgOy1ijCUPgnWsu6q0QgS+tKi7macfd8quIQtsovyF8DhqMNpMr9vrmmD
p4G8Yu+MPdnTEChE9AvKwsWGN6KsJcTqRdmfemUhR5V3fJTkNGnHhlg/dFvDn40D
XphVrxaVbv7jmRKr9ez59cn0aVOszpJsGoU7gmPJ/KxQnMrL76YnrADkqfJdOjj2
aGQdxGSyCRxVIxjxRoY6aPtQFmPMlttkfLmRKiwS382P88aKXVvjfo1II32Pf2IL
WRm9/497V9to84g9XNif6jFkNJLNIB+Rd0LDeSeSZqN8ar2/WJHKmyL+kwyXyBIP
h1SYgtGuq7MFakAf9hcyTr84uJHezyQjvwVRG38uvYIGIYPB+btSbse7XEF4xPdO
FdAhv4RyYP1dZI5C5zeU08IF7a1a3443oqEq1LOVBowxh8eLqeaKgzRZ//M6v4dn
p+IvEDZuFMmnHo/AY65QTvxgbdGyBjAH5EZ/BKyHmvVHatOSt0+xXnd7htXR/i3b
PAaMdQlARojKL1uwfQUFWuZd98j8gE3fE+dNltj8oAtEQ/lCqNqTgN2cAZk81Eaq
kl6sC75/pG+eT2PfqU55bobd5oe9zXCV2G7HMAI2zgaKOHQ9wOdMV1etJVnWf0Ta
xbzhyFF1kcDz3WmisQSxwRZbJPXtr98qbwOzAQAeipvazq9pZ8YYTh19H33R+lfc
M6i+0xh6Y7apl/WFUTkTA0Awg/k1trRVds57ygJfJVtCld9Va0Ts95adq5d+yKuv
w9RhCHL28Rl8mU3o1D619kN772Hlbjw4p1nWcqrW06r5f+mBFFkVzZ8P4ynB+4XO
jgXJ84aR54RhM+jhI0A0134zuHDJVoh4N50AO1nq4LBBYsonxa0Cq5+nhcoslhNr
/tWMz4SUK9Jw2DkSsFgU8U4TEuOpBjN9QjOaKK8HoviTiOa/Z6JRHOulHcK/Qg4i
yR8AvddVRbGEPZY1JscGD0AY6nHjDsXMeV6jjER89L2xoc3ZTj15qL7NqGpN0Vpa
CVyyLMiwLGiKbfTGCjxzs8tnk1NnEmXouhpiC/TJ64HIKcvXywzCaZD0Nu5XRdpd
g/UyyszJSwd2RVKN4hF3WfMaZ5ov9c5tDzWePE0GFaAJVcP6n8jK8zeobyUlqsUs
bf2P2uxkaFmBR2Iw1AC8H4bbDmhy9Rdmy4VDmSOr2qsSVoYVUigp9xUQO7HbcsbA
caRoOu2jZI+DdELfH2PBtiEhRZjGubTDGXdK9//lwu1uQWgMCsywMyzLHcBlVUu0
rbKjgpqACDEwczLZgQpvCtjsNl+OFDfFLT+aOm7aS/BvSBOWyRam+2qrY+Bsjn72
rR1hOnNuZWZyTMAglBNF0kewMlumZhJgRm0IjrCKEO4xTZt1CtFiIzFyaH7Zoxz8
W0Ax49dL98qSy/2WU2kYsKGYtavR/4YeP/0iAlEX+bwP0Jbo7LReJnmi0PvxGVPl
NPfqx5eH63f4rgsh2uByP+GGDh/lqUJiWQGX6eZLqT80dXGr4XeN9h/uOqcBtNTA
MtJIybijhux80zA4KDCgUwjEHWiS8voPof/jgBgddr4UqD3kNb2G/svy/uWzSeaU
9pTJgAS4CG7e6rgzWMe8U4X2PszO1Wx2TCoSGdvYQXCZjM4jcX/myPm+oJQx7XdV
9Gcr9XE4ImraIf+hKkbNsohBBMkUcCFwwk9iFan9aJnu9s7F09j7Fxl8dXKxFQtS
l0vK8yeHFQptmWqYYhnv7XmKfiwXmEFBhjfzBrCcvPe+1r/Od0HoCg+YDZCUJ+5M
DZ9eusN5q8lRFf+fFBENCQZHXMOmcxSNNYAXIV88HU9+z5to+xXLk2grSC8BPTGz
WQEar+QbMKdjD0jtvVBPCtjR8CE2YzexsUjzyyrhGpfq2lwu9fhKhXztWZUBk6DK
l0D196QmQjbG3jQg/LZpPVFwtoH5Rjib5qZZTit+2WBqb7BtMOdFxO284eTJ3xDo
SCgJSB6xZnpmMIt0PPeOSV6ry7wawjA5Aavvl4Eu/RkB53Qmdkh7IUQd4vABWgEI
i2Ur/6rn3Lm9NGNWgBM7oI+bdgshlVD+V2g8iKvxch+IyRxkX1XOaDKKlt8O1Tq3
fak7311H85PoL8wMwQRFA0JAXti67f9mtYqfy8k+RPKao42lBIErTuRAARV8YFBl
4UcJUb/bRwk/5RocatBeQyC6DNSIU10Fw1hMcHbHkFnIy0ZcpQJtlLxrL+Cwf3t7
7IG8VkdPbqDxvyQIxwy7c7DI7+H0G42PX7xuT6u46kwqHO/uxMcasaqaQasahiHl
PFkKosZq+3BrcvdckYUGIvniOOvGZ7gxIqhqAgT9o8ffeanNdl4k68/mUbyD2jn4
McCm2rp6LNsYOp1a4PNmCfAjRVHAhrCNTgBh2HVihUMUvg6AJc5FW0F275ppIUAa
IS8JageJU+kVdsccSrEg4te/zC0nhb0aKXyvum5I6rIV0fBt9dFgbb3qS7MXTT3p
c9VjWAC+4Rjq8idT/BVaaqXs+wGnvEWrb3bGBr8pWxgqm157DcVPKw3wrvD4bv3i
j4rstAfKHcx2wZ5RpwwEQ5pM3ft4mw5hzUIJR4edmbQ/dTlt6a1kF5Qlqni2DFDm
f2I2HnySixYBxKWD2nqbp+ig0ANouMSMKZhOXrygKKXHuWp72m+mVirh/B8Jsj0I
aDnOckW2vhsW4hv/6KWZ61UB6T8DAGwJufAu9/33aKTw5azpJHY11TsM74WUBza6
Q3ZI6SStrQJFXKkZ1ibiO2BdWvtP7vebfBM8ct9mj9K6rF1m8IKPqEG0UkxaXMLv
7RB/yeQBoA9Dr162XeL+YrQX9st+6dbNYo/YXHPC9wPlCOMW9s707f1bA+r20es/
n2nL8ZBRI3qcJb0WLosiQLWcG7/m2Y797qs8FZKCa98CF1W/XAuop5Xx6HZeZB10
EeIHGRumhGQ+Fa3+7yVj308ushuxwExVTzNLGBJg/C9e19vS9+m6dWFY2dAqN1o1
McQN51GvZiIB7JTDB0icgD5c553vpA/sxclaLJ3Aa5lL8apIePIGOwVW9OcZR9T3
Pqwvx8junV13ffWBYPj9wGkN2vTGai30/UQWI8MUSDev9aEqUrq0cO0UibPJfxDc
13s3H7MzBpL57LZKDAr6vK7nWu6UWLHB+oOyZnv1hrk45GADAFnd7TNgl1Ia9cXq
wmf9Z0YkAeVXwAX6cuGpdaZspBnDONjODPQ+iFiQdDlOj10KNKEqBBSkj+LBgGDN
nCsLwN6lln6w4evdrgJ+8t/VpqhELY0qzuY6Ux3PWhPYA1pvvQWFGfrjvyfA5vs9
/ufyzIM2LObDXglUePlchkeKxIQpJ1pgxxBYQmljreY68yU5Wf1no+MqY734ppWN
YR/EJxY6cdDMkSPT+PtjPkKrqobNe3JsgoquxLTXqSJjCzkJ6DdMbpK/9LLfBd00
lc2/HS2Vrmx38OVlW4w2C/2pRkP0N1FQ22GSkQ6EXkakFN7xLqdrfLlS4msVbUHb
PXpMLlweKgfMS+8JzJ9p0SWah7EtHTm0utJ1qiBYJxNbtoA36nbnD4yit7rc/otb
xlBDA/sQ0WzJsZu3ZHsHNEThDapgscovUYmmCG1ptChCImtqU8kNKaZV/0sUfi81
zoA4WLmLlf1KT2/IZBFbhrv2VmkRk5p8wiCRLKqcI52ZVDCbmzP1vE4P2DszJFu0
bcHIwefby+UY1CuvcjUfx2a9dMKijvJhZnihou+2fKmd+JXx0YnmNt3TtrOKMmVo
D/HkYT0jgVtAPnujUesZvAjLzw0+CxaCwnIXJ6puPtgtTSepWZpVI/P6n/yKmSh4
2pbVQqS4jP8wtYU8FsEEm4XJguCdMzcEsfmSBk1VstaMNxB8BqxKs8r2Iqan2kPZ
CZdMLA6OtnElg0AB5TlKia5gRSSp5zKuOqW8ERuC6eKPlrlqKD9uj6SafTGYvqnV
SA+5Bbx8LrozpoQDNtkBWDCwJoUl2Zi+gazR3zwPtIx305K7Gz2TVLGoGg1jZFI1
WwfFXVzwXZBGHJVEBhCaxjKZNCZbuF5nvD2g/KXE3hQOV4SarMMktep24zPeVW1G
ZZCQT7eH95SeUOzTpucRDKiIjunzFpiD7wzz6sM5MVSH5vgxy6xBUMezv7BzOK9X
awI3VlfBvX8+xo50tKa82dgJZfCb76JKxeXUzWs6fg0WfdpdIkF0eJegIhbA7cvz
rI6lP6xCVCuPwQbG/somVL9chH1QMkEyTXAHre+3C75tKkYpBMZQauG7z6Qb8zC7
OfepyEE6SgqGim/a634cpBZU+d4jBIQJJ/ShJRMiM+p0ewT1NUnZ6uBlzx0IXKGc
2EIRO9WRAB9rcuMpZC1jawhxoDYF6d268wS2GMdw0bbrKY+shy2VGlDhRT61K1oS
BiGJCuOfTc4EfeaYvga1jbNDR9Ya+HOfqrtkQGeR8uL7BUg+4Va6OdifdG7VappO
M6O0AZxfHdBTp7oNCu2p6Mx7fXXQaWjvDMAfQMcE6CaEytPdb1n/KkX5p5v0iOaV
4Sgwl4HHzu2mRkSH2IUMWIWnQgXcG79tDBAz6kDAQ8oYp7ALnB1xLXrW5puzsDt3
htNDFx1RDlBx6bzgRzKcZTAx/TiJKXEPsZH7v2kRUMNhfzjAdHfpqsN06fK1vxeY
rAsjtkfyjXvjeW75hbIwRhZteZqMk5tBvT/njnuB4lyqo6WS2151VTZ3lIUuf8LD
Snsnc0URXaQXbGKHlHBsJsQZW7zQEg9JxSMpsS/DiSLQ6e77DN456oA7SaGq+qHZ
R2AgliphGcj7EpqWA9CPf7MFDJnudaM/uXMbWJhrje+twimNfk6dhyD70B3DxODJ
t/fMuZ52KIROtZUBAu6y/s2aBjrWD9UdHYap5voZntIY7Y2GEYTiTb0RqKr1qhN1
u67HXwzFxX4qua5dFrISbWwrOkHmipB18VSQNkbmJGaoLZ5rJb2y6ZtQTGk5yYHv
LOivTtj/e1l3RbG5lgdS2R+dwAYEP7wZJN7AWDPwOQoIHki78oZGgnKkgTb+cvLV
dQDxos6BcAXIMG8fRyviWDvAVOzs0g8FBN3w5U6eS1PQ4QOomS3SBsS1C8BrgoDS
0GZCs1ZGHxuwA3942IsY4J7cV3M7U+9dBZwxfUas4vAddrdtA9BHvHOPc9u+AtiS
l/5Yi+h6iqftg/TB861SCvVJM1M6OpPwlSTL8jXeeBXyfE5Jl9FGFuyDcMiThK0k
QFZho0sCa1z0jMENJB1ERdfBpPQB0SfbsFWL8TaYv9Qb2t3NVWrAnPhCdyZQypA5
IV7hrwvroaz2W6twiDHD2ffDHAMBi33P7EIEaNkOdh0dCT3D8/bjQfjE2AeYbvar
wj5N0l6XWj5NksdhCzGGh3zq/h2UtlrHvyCTAeUcIkB9RuuEwLsXxuMSYcRUyn3Y
je9TMw9cNlLlHu/UCpdfotcAc1T6k1ogto5rg/BYSqyzC/WUZm0R9T8KJrGJoGpH
v24F/z0QYsL1qDgaoKJSobdAQdyhfKCfveCvKggNUCH6AYHbog3//GqhFg2XHyAa
hrdQQSg+/NbRc82hrbxB0Z3lvjfpnyGpmVrfsOJpghMobztk+N7zsEQovChRDvFo
wC6V84wb8ZscqLMjSMcpiIXuAdPX4tl9JP94H7h2spzBDawTD+2dpyK4lmIPlRqo
I1tUgtRf1rAbTFFRc33gDRpHh8VvcY9fHQ1Ire5L66o6a5QqBDGczZQWLNkQYkbQ
arMEf6IJ8a/MVPw6DLcDgWJjyXEKj3w/c+ht0Mi3AWf/ZsTvgEBFU4iJG/C12YlS
RElwAQIgkz5N7djGV3OFCKaDlm9fH5to1Wbe2M34h8WOG+dFghLkUAdy9TYbP60E
NN/o2WQX2p9f4rwpmugfxCchKEAjh6Xv4ZuSPlAT026VT1UBw47x7xEsAOc7aXYo
EEvRcXG8Jojojtw0o14tzfydoxNaD0JvyPGCUB/3i806nouqgsWso/pxNcOzK3wB
vAfVnHetNuS6Nc9B0YKvBbnDxkT/RVb4Tx4wvdIqT6sFmhyzm7Imgx7BgQ2Oqf/J
ov/MCfMDQtDm2C/Evmys+cOAwP0iylk5wWXqhe3hKQuDRVi/yY3niJtQLf9fM2X9
HPM49cBCDlW9NdhgO3xZOgmtnx20E33c/W8uhT6U0EWTjsOUXU3Rnt3IeBioUTZN
7OnKB4NR71JjDLuWN/DIo77psEIye1aEYGiraUX0SqCLisMOktfS6CLnxT7sGxct
rnbv2tcEUaakhI4xHpGYX0eYwgDR0AYvS0pW2n6biXXqAucGcY9WKte6KGltJ01G
KgvhWUGnjJfqtNy9f9Sj27QEN03odpgvQiaYPcGPfT4pSpSpyf6hEg3zrsufFOGL
KafCfxpcG1EH1maeqKTDKVDjnYf9bYcA8gZbtDt5jL7rTuRMfD1dnudygzMEjrYN
Ky5979Dg4PKFizOic1Ed6487BYJDWqXESMxPfdP+L1g2D3jGDf3/jGYghfkEotV3
axNDYWOnQ4mZ73KjrG3+tkFF7bzbJJiYuWq/bb2ljTRyR1yoMgPW+arn1KLpLp5/
BgfOcRoLEjDKCUIHhCa0NIEmXxJRx3CnsEtT69fnABvWgvdM+ESFAELcMZWs9ccq
MSyNjxCLjmYBchxvpLNrZiEY4H0otU1+zqqwdnbouBxUoTMKWT/UFyxckgzSIu0N
Z1sO8WWcX7QtMNDMO+7zmQMbRByO7icYSybza6KJ7vzprM4eZkmRIPcuJIrEcxba
QzZ3cmWKn32m3ln7Qntnii1lFwQiqHbRIho7O/1JuZ7HnJwlgsD0CheIM5t7EY0O
7bkde+37iiZlwYtt+GyvAZhDzix1/yd0z0laqOYYqcrBw1RoLv/bPxympPmsYoQX
KZtqvVVdfZXUCJFZGLVD7cvG5EC9TvI5pAdQPJE8B9JcU6XSJFaIY4Hc6kn8BYDI
BCwBBCEIEPDXHPsoNEP+Zti3jG6G73SQGz1nuKrUjChl1h324cvOWW1I8397zUs9
Z0zGlhnqPYFPzoOuBdvwqM50iRV26Nw6lK9Af7lkXi2UCoXBwLwtd2LXGlARf18c
6RKo2jt/XOqxjdIPsMUPkt3/SUgbZ53XlEpTDarT/FQSVjJW1W0Cc4afGtdVw0cO
PtNsppUk7yuiYitpRWlkiaOSgIJEdx3AdNh9Q4DIGw2iaaTSul77EKS/qed+AXMs
vEtkghspla0gPFi8ezYPaRZax6ubOIzcUJQtD/CiFzl0eBGVSiwWWj1lbeC1CwWN
mI3RnrF9dyXY6Cn9Nik+KjBV/OgPOewTUtXeD3tQVv2hBCJK/ynI1lMD9iasu6PU
cgYHTgdo+xlu9qj9F2eyegoBbk6BdWzmtSCa0q3oMuRyDD7kjguY0yEOIMsx0nFh
cd2S9UjcNJ6yQljGgzkKZIm6HCeWkKpp56vTllUWs4WiKghKppNR+nmqth6wZqRb
8xMGYcZ546PLI//GuUSH9rWwE1jVWT2UmAXxyjc9ds9tg5+JSeJLBlp4hTU788dV
qSEpaxwZTc2rpYxGhi2JkxG81xQtQ6h9pxg3cLF55hxEKoqBUvc203oXvXqrWiy2
1X9qBf3adE1Dyw9efP4ovUhqW+9ClZ9DMzA69pmfhUyvDFm8P+owSWrbmIqopyXf
SDsIzXqRAPrV2sLQy0qJU5lJcyFmA0YlF4UC3brnjxnaz7j7RTArPEVqGBzw9Vu4
R23m+y7H/OK7FNcMMZFyAN4NvFv7uIL6on/ZhETJDCyfuMlk4PRGjEs04SrJg/+C
EGPdgucM1Z4+/dgcRUleCVaJGG13+aHukZd/FGVlHP2mmVTBUBAyqjqOX7u7TVjn
sOYF/bcMADRxluDC4a6XUt+GfQsfls4jlVC2QU8qrNXg37oMK7FvTM97g6jYZtQR
QAeXy1P85JB8w3KWreAKd+JZ8nDX8UogL9h8DXuR99FJfCvyH5pWuD2fCYySGz3U
f94yB5dZxGc1kyxwdBvto61vvuw2CgdynO1slNbGX19eKBGh4bZqmqB/IMbzvq9Z
xalYv1XHcV7CuX6fMgk7DCYX2fDcvYeQZClKK009mdjq0KXM/KxrN+5OBTWdLVG6
XSpxyHc2LzwyaZqHPQR4jMYxjPGbUHLIxn1BGM0RWguvkBvayPJ5k2a/jVSH3KH6
hoZaLt6LQ/HEmRSuCMtO2RVDbXQWYVX9oTt7/zeNMwyyVPVddS62DEInyxLqHd3N
cuCxS++7Tb/OuAEzBL4DJoj0m3FKiCSCU7zMlp6l+5oxJXJTAgHyX5dTRS7Q8V/u
TG4HsWgrrGMWQXj2XOnauLDl4UufWIuCR6ir0SJf8ywftYD/4Fc49oIvVUfNqFQa
SYh4rwpQcSdrY7WWGkTr+WAt58X2yIZPPSzYpi3yLoejWvim/f3NJXyWRt9lSJJ4
+4lbf5fAnGPO4U31chZuJpMy6jh3GBjHJ8R/lo8bHWRcnSF/pPlQQGMISYKkqtF6
jb3tb+D4q+kXklAihw12ccx9TJzMguTvbvwZ1Xpf2CkjQVuMuBlwlA4MA88O/62z
oXTIqbGKTdlBIfdjZHwJHm8yVNNcHaws9qNP8BCeJz9bH4nnuuogVSW8DfbgCj9U
2Od6mCkiFIirqv9D1OkAGXTvWNqsyO9kPF9K9t92k9d93X8IaoK1LFORiyWqfVFr
yN9eOw6su6xlcdavCdd4pSRj8jGjBaZgxcAZx34EvLJhm6zrVhOHRtd7EJG7CZxu
TnD+QyroAbs3Zc4w3se8qzjyolbvgyH/UTHpcDPTcWKCQS+MsKS8jp6Vd2Lfi4K4
E7wzqJgBmt1cenSL4v3zx8BRWtMqM40feajqvA+DpiZhYu4bqkWG6eWdO4Uw4vnd
6VE4SaXtWHK+UBdDx3+oMh3Vy9o30+n2jm8LhDxJuwjynDXDYkee2q/XuBMT2eP7
y/GGXYmNveb5D1m+ozwk8RCwj33KTrALbrnJRL16y/dInv4ioVaqgvr7vvGL9EJL
y1y+8ca+NZcfXyRRw8r6oTGbsFhE65kBlljpcbpD23/mR8y2oibVB42/ZN+ix3Q/
2icJcUdj1MNqsZT27OqVAGeDr0N/VffWksDzm3P7bfZcJDqnIUuNH/s4qcRhxiV3
XgzNk8dvfJZ48zpFv0aL6hsTGzUoBgM6VI9GNf3/BJLf8MfwsEpSGq0w2R8xoQYv
vjyypJj6tX+WavmWD6Z2ZiORBCe82Mr/7uX129eQltlMSQmyni6p+hi/CwSZXw6v
nVrgX8tg6kGsq2Z6dW7uv7tF1TGrUIBtZN59k34VK+khXYW0nV+nsM9HfMkgvDaG
nxwreetTRwfP5L526k7iHHYwT7ccA9n7l9VSLmhEqXHoxHgtYjn2y9/CxXsKFRRf
1aw3suuuFZKwOpcDJUbF1gkJpQ1BmCQw2W1N/NLvFKPYNrtVznNkWzfiKASCiIUE
RS5ymjgShwsnRFmbYw2Qks5vJ+dtPHA+Forgkbf4u25LMJn04rfq6HxZLztrx0bq
e4YeDWQMslvMQ3raGBY6LDh0jC0zGDz06naBhsxIG0GsXhHCBpnRlvalx33IFr2O
`pragma protect end_protected

`endif // `ifndef _VSL_SB_REPORT_SV_


