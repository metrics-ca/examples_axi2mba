//----------------------------------------------------------------------
/**
 * @file vf_addr_rand.sv
 * @brief Defines VF address randomize class.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_ADDR_RAND_SV_
`define _VF_ADDR_RAND_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
cvmHWdSr1hG90b1vjMqAV78HB5h1YpiZZwudD8Xiit0JutdG7ZeB4+Ghyqs8DMwX
HLO/UBWLXry405wOYeFldK+bhoNhWNrLCvZBg15YVzZwTdOFHm729ET/0uPo5gZn
OMgAfTb8HWtc+4RSOGIezz7UZY3m3ZYsJFrJGkTDCjcDEe6oNZdgKScgGPFEsEzq
7/auuMDzSbPVsnwopgjc+DeKzQ1VCqUD2FbedVvI7jpjTe/y+nKfENOo7oLJJlza
HrgOUD1me0QqKFUFcv47JhL7X90hCoBkhHewGPwrqkd/wMpOHJ68ri2ZsChNXe7h
WeF7vcd7+jHvBk6G7Vm6AQ==
`pragma protect data_block
c/lf4t7a3168HMxvHZTOihN92C21OmfBdYSQ1d6ICjdkhpNms06olHUVHH3klgm/
mkfHzax/Kikipi0tneZlIs4sKQw+QEoHRVrDSSW7Ui2X3jI/ZGbPcrN1m5ZlcGuK
T1LK8a4RWMJzdHihLG+gpgkkiZykOTOPeckOPWFd7WgSJD/lLVj/IyZm8QYvkY1T
FOrdu25d081GrWjjpi2AzN3yn2/AS8jl0O0Mn9Yb5gaFHTIMMGGTcd3x0B1JpHSs
VtBEV8V4LBSkVYITmKmUTydhrc3oV6T3S66wKX54lHXdpenfRZp3nz5WZWQZv9Qa
rVbfvjfq4u/KwQ29LRUtY/Mc44Z2xyudRAgouKwNt/PkU7XCVETfPzZGKpgWG5iK
FkuJ4bCgYJAr14CTwUvCKaWeS4FKdfVZKdddqfrXHItQ9VgmWTKeplvrPn7tT+ke
Gy1Xi2w5T014cyJYA2sSnaOhzaJPOMp6PzNR1KOaEGmV3mJnlJtf0BhX3W4kBJI4
HCqdivu4ld5gtBvdSaeYgoHhnrAariiSyJsvBf+FlY6ThqINtji890ndhUGiyYXD
7PodRc0Bkv3P/Gc7ZAvgFYzKwQYH+54166+446OvBVWa36S0b+px2cEr0IhW3G6M
u2m0S1pwn7EIh1QqzHYjRC2WvVE4QimhKNfb6EbXiAEUMRzX5g0BUjdMusZyKK6H
+DTPBGRdLdDu8xIU0TjtUfEXdJJQoTJ0VigpzU4dYmTgQD/HF9U4t1ZlsNs2l8lm
8ToUggDHzzsXZvhYUDtwfFxJm37Kwrto4gAuvu98vh2Dr2vyWQYrxpdK8tGKyIFf
bfLrMNtFa08qowWdhElT+h/kzNYhcPZXtm7rLTwIg7wI5/baAuIJNY+FgTgRS8xl
kzkeeT9QcgvNjilD77af1luncODSrLoLHE7ERfBzuYzl9peCSFhBH8WP+JE9vu1+
gBVd6qge0jWTIOGSd/FZsGtg3BHSCII108dJsON0z8jpbusGCJAKtgepuwtVQxoc
4BMBWAW7Ojf9/dfL1NakA3IxcU6NjXtBmcauo4oJJP0uhovtfS0w+Kpp4hMPx5Wx
xlON3Vw2S1Ta+QaAZCZTJV8SEHTr+a8Aqy0PNK7ldrVXgBt7Won/Jvm+mqRfb2IL
X6qJ+nPujygyxFI+QNFS/Mw0QzVs4+TPMrJvgQMnFJpoqOWhOlI6D8hM7vxSf8qz
kgLtxhDOMiJ589XMdTmPsraEVFI8hMZbjnKMuO//02MQ9cFFHltWgDoBFS9OHvi6
fmrUjpseW63AtOPsboOGjrws+xtkCdL4JZYZhQfRWi0wJ714vAgHcqQy4shzCIvE
pHWdZBIv1yHKVK/3KHJpxBCbcbToaXgBbcCzkwWpAwmogKncS76V4IpjlS/P4PO9
+0dEazRpAfppFWO/gNEeFPZ9jgCBPUS5h9sSdBZee+TtgbiT8q1I9ZE/SJC0jRPG
KABdq+UhDbe7EJqy/XMbSn50/gPgc+NeZ2qzAbfM/hTUYbGIs5id/zA9Wyxn6gt7
K5TYdfMMW86qDzo8ufA7TSu4FjFpb/e9DY+ZzJ+1X3Jv9uHjnsn3vxxZ4HXgxvBT
uO/6YpAuWtaO4LjSDlD/65EXJpCA99rlBfgRDz8Qp4LHqPVwy/TsIoZU9eIP/Mfb
LH7DDASUab2rdkLZXAbETbLSN7FnlGKAuh+HVAL5Bf+J0OyM717mgI2dzsP01tw9
XXSPNJ79iJehJuGXbBAZ3damjNhH1YmM5r4aS1FmaVcHSvecW7kmrgHZGl2/N3kJ
orwo74eQAO2dv4RITfIFATxhef8+HI/28s1O1jS01ulJzY/u5mv2N2eDhoJ/7g9/
C+bclXSo6udLwsmhuYrAEIP7/XHCgP9TPoagWx+EHgUhzAdW4dCODxz2ERucBohI
c2+D0PgZKmy3sJNJ5Jk8qH+AvZKrg3lTMPiIN/Z7r8sGc5xFu4t7AhdHihxY2Uso
pdFF2wNhKR33c/cOiT79UNJta2GsLhO2jI+2Un6qFvU6X0fNU1hQxr8CURxMMcDp
PmaExrcINFSORqokMFRIeSeJaLh7SeRmnJ0GgS3dbsgaBzc2JeJevHmliIY7pvG0
kEOCfyj5P34xnEHyi8A/W5mLnnl1vg4ZiN838aK2rHy/HuVh5fSEMpCWYvUiYhsd
V4p7jzX6acb7SVtCffqYkcOmuD7WOjgpycpLXsUjV60s2nUbkbStk2gbi7/GMRyE
Og1Nf8QMkFseJ9SJoTYQNcYV31cU1NM+qXADAk1z+d68kVSiC3WBE51oX3g22Mbm
Xn09pA3PJoMfyru2UxmTX/dIClEaax5SZSopfLUlrMH8prkx3Fyvlq/AZstRtmUD
GFjEgDiKC8CkAObd4zA2eQk8LzCtI1lbRZ5JkXr5uuV6LOYkoxmPepqUZwipKYQS
3z1YHLKCKQgkmucIFz+jUF7jfGpp5OQRZeKpc18C7ukw+WRCd6XvVLesKd9k2XL2
iSXilhT7j1VnGVnP+FowI9GAQhviW5rnIV1SoUfXvfyrB94OlJmnhPsY8y0Uzt+l
2+WU/KZ/EC8ORqa3wscf69Th0V/oOIp+WIFgFNZfiZjhgujiojL/2HRROb+Uz5Hd
GpUFer+TrYUO/EU320r679B4wLbgy8tWl1UzRl8UxAQbAXcXn+w2XKmwMrimg+dZ
kSdwOu3MOndg9VyLawws5Ij8Uux45+14+GU1fSgJowhGT0iaSCSOxiiwBdMBNmGE
NW2FGecFmxO0/WxHEZe3/jsWcGNhq67pDnLHl0CE6EE1ArA/1ah5lN6EZvTX6mk2
GQj4xbB5rBdESwdjaEeHbh9IZEVoQVYKziZQi+u56/JDULv+0ce+rFDvldyFH2vL
mU+rLIo1sVT85YjLidCN/Sgl3ulU2QXd7mvcq+V6ttH/Ob9iGBRN/v0pHF+yJEn/
teBP1lSK3tdlu6qTCeNt7r7YZZ+0lMD3hLRrO+URdLIixi6wAR/6rneMvzFUA8G+
4fxA3Ok0ZhGrM6XXzmVNHWeP3vPgbysz3x2yRHADIufuQrm/Qq0WpP//Qb4QscFe
nEB8ay/sN9pLR8KDizYlZoZZO39xkSQUof/jJ9pIf5vlhZfXy/sMZWZcfGb4jd5j
oWDNNbDubrCBK7qtY9lfnA1V9XxolqXMGaoL8lKZg3g4JHHkxyEV3Q52SDWL+gQF
mk4aIN94PtotNLFWfkNPLyjpiLesoLPK8KrKUIi2iXc1bHtIaNm5WARPHThNhcjj
xcCsG7OolYC3GHk0M0q2CviKGgTvOZCEb/enHyKJ1SDkwTZGJ/m8fylSrdgrpF9A
lpNI/DYjRdRFhbfztnI9wUp755GnpDqthLFU3lUcqFgznG8Buyy3MAxYUBxn8fOf
cQ5EQv3+Bmm0KC35lDRGS1yog2vbuXKQBLmPiOLg7JqeAHRRPt4LmKkbQrTTi3FQ
ms6rN5xtIihV8LfJiIUD0yXyyHCpNpc0GCGlva6Nk28j7GRhAdgr95DaQSyg5qY2
AF09kGrwRTeBcv6uL5+kI9kDKCgRLqqULmdHyYfdwhm6ownUzjK9GgeSipmpwWRB
VzfG1VoO5Rxri2zxQ5QhoaowzqBhc0yFH1RjsEa1HD495Htl6yj8ikDIX8VAQ5gL
zBeo9zUAHQ2vOaie/Cs6C7xfGBvwuC4Vm3lw2H/hjDDYgKlOOr6rsfFRSRa7GY4h
k6G7gjc0Jz3HhJkJmKVePzdlVNcLkP0XgIDgtUgzKH8zbTh5pd3mqaY3cxoPYgcX
yrisa6HXGzXlPiK9irCOkwZJmqB2OVCltSD/Kajt+uBUdfp3xbeKfBz95V5C5joB
yBHKoNvHnm6ng8A5B5Qb/yp2pSMz7ePObKhLZygKap5suqtOIx2TNFqxRpIq6cOB
OH5XD/xyQ4Vu/FN0yFnQ9G02fv9qSa6ByMoi86sYNtLTd+ppdXz6Vm/VlFQM4lVj
0L1ygKJAm0WNjvF6HoTp0KD8LgH97ogqJfKaYocH/l6mWHmxd0JMkbbW9Wj0K1as
gAq1SkYJF9SJYiM4WsQd806uGwjRvoJoEZl6TLVsXk83tLogpNTzo9eSQryeTKis
88X0NOZA4q2RX0qqXwUUk34RB46KpeIKkeV1mGkiM77Pb+LN+8TVDP76f4PShdzh
B+bm1xCrsOlrO0cJJlkyPzHGJ+qAkzpEqKHUfGVqAhXohx8/7eynvtU23C8tS6Cu
zXVhtfxgOuA4GVmVehH1AcLeOxJ5BgBkVKusngNCno+dAN9639PP/hoEIFIsOZVe
q+kRQJ8EIctKz2qOMrozOvIKUhOWKcwruCRqLNYFes4HbPNhr/jp80wf5A78Tf+h
+8HybI5dck4fSm56G/X25rrUmnHprs8KQSvQ71F3GpDgWDhgSBbgNP/dgHby+WO4
80jRZg1SKlcAuSb1YRKcnY0wBxr3FHGUY2qYY6Fj/VQx178I/YlR5BDQ+eweuMhq
OzAP/Zv3HW1zGMlqqevbZJ739P4/8kYaC6uDS4LH8E4qJtc+D83LpU4CJgHNLtpm
1x2qiTwN7ZmmqS43PZNcQ3Q0nd69ydR433HduwEAmczCTZYPivn4qzI1LIm7Eksk
0ujzsMUNILGia+ISky/uNWpiALY4+v2RkfgYD+D6tTdTo5Y+wo2d++m9XZA+wh3P
/Xs2YQm26/hymhUmySOKRNwYLsj+gbzhDv99hYh1DVrV1xUB9yuoX8hwnHIkJFpY
CP7LQaX285nqTRxg/FzyGChNCYykZbP+fn6ukbl9XmWraZCIcgZH5tXA6p0Gifvo
lx01Rfs3zoVEIvMzg571Z1S+w8xRmvjivLF5VC2phZKx6CRZfXsHj7w9atsLiOVp
fa30c7xcu8PtI3B3zwgHZjNcm3SboQZjHszHP4PXLcSONWLpw9rk0comKiQLacnn
XKPuvUyWTmy1jPz/AvASKASeGc6XO15PAgctUbgL7OEwwvKvraFPMpeH9/ExapU5
YbEpOU++TVm2o8uFfzhN/8862glvDdQEGkLfVqFNZHA+7sK56NZPUSK4ej/2TSiq
56FkQabMVAP9GBhhPkG3P5R5Oe+XNUdDRCqUEfKMYnSN4x+iZOCPV6KuVrP8OvFN
euTkI5Xsu9CYUHoK3R0SW/WaETpdEkFGam9t7YjoVevBU96PvFJkeGDGyVOouBPp
5A+ayUZhHA8wH1XaFAFPSyPLoyO/+U4Id8Sk04zHevPXRsA1DDdrSY/GEyXovuIc
P9/C3Dp/dfxT2Dio6KPKACse6kYSbK9sUXdGL8uBg0leYFW/PiKEjX9z1vtDPGrz
H9GFPIVVTH5bUAhORTKtpkikxxTS4Bul2awskmnaxAC0i4jyvu4OmPWhb9j9lSQR
rqgKIpeYUhAJIpDOoNqb7xaYeRN4n8Zqnym+W9pFRcu5OTUSCMw5OtG+X8WMFngc
smYIk9EXLm6GpjoSE2ZsQ6ZyzKvhhC2W6JRscTcG7spEk9sA55eiebBxAIuxdi2G
2rA31n/B+8krd+HVjT/Fmv0oWdT43d8BHuHazMbfd7LfOeArzNl4tff26uiN9bcs
kwTJ1IyiycdxsWV4MFEHKAlC35U79ScICskHyORHk+ty2gPY9TEZIVzZIoo7sy5H
0O9sENOs4dWuB1HZDHgyJWRa7UJcMqWOG1litHcQs9jsT2ku8c2PqJI/TZB9BeOo
F22ndd6fvRR62Iw2Fs+IxwYTFRtsYz0pkJ/nCdQKhFtkTI/pi8YHVefdV5EYUi8o
VvznqQ/+BaWUDwen9TwaEJL6UJkV6IV646FSSc2NthbWwrICe9saDIHaEAiWiJKp
NaLecLOFZvYN2hhZEhVKaIL/9MIldqvXACWPZDHedzW81Um7wRbCXZu7DxNeIigF
btY0OftS77J3ht63nlCooSFfQslp9fxMChB+gCsqb9R/p2mEgFIqLQ/n8YLV6DBp
9FyQKld3W/0G74sw0GhHPyVF2c8BnaSzWGT1d2IcwUOsVx8B+vGYVSxRUrUZ09JY
VlhdYR9FZoxiNuUxNVtvKPUg4ql+tZIZ5kMVsdC/DeDQObGhtZIjP2aAXtab0UXA
NW9USrVGO6jDE6SdQIP60n4fg922pgJwF7O6MpMrxgPOMyuGU452piFy1K+6+qrA
5Gi5v6PVDZAAHYAkNW6ZM7xsn//+n6NXzf3iFE8sdleTzG1VI6q9FSfQIPjUccN6
8A9JqCyn6umk7QDM9Lh+NnpH87xvvdSiPXOvZX0geKbnSm6Ua0/Cf8SlEiee04Eq
501yXL8sxEV3QD3HgV9R284mvZyhm3mIX9FHP7DRxhHpU+6laCj1gfwP5wh3jfi6
PGW3saPfaMECCvACWCWKpDaTfCZ61H/Yjg0wxWsleYxuukW/fiBUFhqQRHfsxU+7
P2C8clQZLEcq8YR3UfDzwxHZTomxF58GeSNk212Z+yhZnbshQ25oxpiKgH0nXyWC
KJVr4ELOSj/G4/a2Ci/jnYPdPRO42kmtktgV3EtNNsHbFJtjUVeRycJmAKkCx/va
SYawVEzfqYdbertaADISznXNv5+Ayb1TBlbuKa0SUEA/7EEdvXvsJ42U+nCmjkX6
HtBEx3yNsPqwX8J2mI9XZRwdBr4ecnzq6uDP9ElVUdnRQv1oxkxkDUBwBMo69xfm
TrDzi6WcNSLwkoZiENl0ExbXmkaJ8kE8wOR1+1Aw5PnOG+bKLnUt8D14DvyLvFt6
EfJaZxYu8KBkQvjjkPupZcihoFZwV5pSXyfkHSzbCGrkKi6fcRYL4h0esK+FHQeE
KxxlaQ56IBR2fEWYdGAbj1C3vvaZRap6duc1b+ZD+qsgVoSkiQpRnMFDGPCEcIWo
kM63rkLg0erthwM3WpnNK0IkPBzaD7fGp0hDf0drD/aXh129o+oWrKMMxxyuvhvJ
XwhIzIFB4SN/bwdtpPG2Hn12QtuyFs13uLK14sbxATKpv7OqaZPm0BnNtnEOxidX
+J/ncan7Qgv5eiXgDqwYFv4cWu/HwXgRi3nDeJ/8cJKKOWPcWyuVMG/4CyEAAXXu
q9Q62xlDO9PS9sHw4BpxY5YpPsTnT5Uw4Z44Dytzd/SSt+Fs+WlkdccA7P98gI/i
RkQKGyIzxdm2T2pbejMuUQMNJOjof9CyULc/4f6SGhR8tt28rJfsx4BAk3X/NoUN
YtarS/SrWr3B/9i3hqVnsbIgMf0X+uMQgeZPXyOtP0y65KNu7UebLbEnLpReUHPu
kjt2SLFuoLFxiEs+hc4qLDmoCalcEMZp8jmGZ5GIlxPmlBao9OLsTrwRy4UgGngx
x3zcDwvQ8cOyN67WgAgHErsGjXBrNhG+1dPtaEO9uQRvkdzzHdyOcV5Odegf/IfY
iayIxUCAWZcGjIsYuRP+K6nf6naXLPBqxpECYPfuUImkUg0G9KCCbPsdHA+nWvGW
UDvGu9tvMvysEAgmgwIlwt+2M2PyAh3aSz/ktrkbIMVd23Q1EkAvlGMNcIrl6any
Ogkh80RMZT2rR6DStPEkxb5I4nUvcjh6X13y4OwwgYy80qg3QHtQqwFXw/P+8jNt
0D7oIQSiJ0Z6Mt39FR06hhVz3EHg6S/9Sl97Qx8XKKsDfsk2XkHahrzWFtGkdiNU
XiBjzgeyrPVF+scPi8aOq7YajFnWwdMN+HV7wfgqw++PeJH1bPuqC0dOir+BfZpg
gsnqsKiee4ovuKUch92pdF5zfaPjEEXjzsaQE0t2Y/wbN0bXnJLY9FuS+2A5wBL7
73wZlT5dJ0WmGS/QTQmuePKp8PTlM9KqwQ8/V+5WGyST3oqU2HcewNlEeGUZpoSY
Vfy7o+p5B9IFpVHOi/cuZTqWZ7e3sOmWjHjw0m3VJaGakVmdVCHYVsS+ft9bRKB4
0cCSaaeNWR4GON56KUo3TKMXniaMGVFVrTuLXBAC/ybfpZ8oN5zFayJrfMD361Va
An7VtB2PF9ylTQsVTl95PecfwHFjKtoqvkZqFfY8y8K3t5yzBdnW9jUyVfZwok2a
kp6GKvsiGpZq6UCcwn597uEzRIeMnrqsaGTeWyaCDrSR5IEK9gccRHa3NCwc81kH
MxQGBbVLxpDh2cQFG6Tm3zYZSsql5tTi0XSFsJBiqJYv1hGxWkbWQEG5R7zkDanz
aBNomx0jCJF77LJ84xKZkm9he1ScvGOKx1G1xuiCJ7WXRnlyu+8Kr/v/aj47eE8a
Y6Lr2ybSYGgukH4NQEtm+VR7G3ksm3OQ86PrjkxzFpTx4Qx2g5ysLqnKStg7y/2z
8kjLCOJd77mEUOfB2fwtw/h3QnMi4LvHTR42yT6GH6fa70hGbbtoOF7FeT3tZZ7f
3YcVxeDEXI9trostHMhBOS1OcnPzBJsYW5n3f2amkdxBXU2LEKdms3tdICLmx0pE
U+FMcXiT0umyRTFMKqkGjRTNDmCmy4Oplz08IGLjsZNfAWXKtR2OmaiqY/yFXcM5
LTMFkN4VAb/6XGraIGk9IfmIKaA4uPGz8pcBvQrQGe0pRHxz6PI9jQyhhyFLqU4M
1u7jbsFqgK4gkFRnKiEDf1VjY08i0TaT5wDVKcKnlWKe04UqXG8uQFZd1VosyglL
4XE3ZDQ4hJnFEGQNO86o6cavEOxyXNf/KX7k8ESxAVwCvdhCsj47jHMwHh11u8zg
viTftEgaWwN6YsJK0rynO4YMPC0JIjrl3LVhu7S8icIDvYDiNgzAEVX9ytC7jFNJ
3uq0HodI4+B4+xrau97tk3LVALNdBdMGAljsut3HQcoDzxmFXvWFobTCoz9rHRv7
yqntemeZUA89yZKKOcNApl/Qjm7jrLGDmiE6EOIGxnnMxva4GCQv4mv41F1gyYc/
O0mIgn8LdSjTAGq0h23egC/lcNu49E2qOB43FzpGlfuEtyJevuMZf8Z2c6mectrx
jjGLaBG785Ur8we9LhgOA/3sQQ9JCy7tmOsi7UvDhgYjfvYwGgzy8alXAlFBfxAO
EmC3ZL3L4aO/5lHwnpF/w7wN7+2KaBWShRNEdDQxyQSDZ7EBT1ibe8Fui1h7hbs9
IDNKMsel2s3socWHdj0oM4DujyAf1bz7t4OJWmvLVzYCCdt9oMReY01h7XbJ1Zen
FTVKluQhsGFN75UnvhqLmHh974Ed2svzld+TEPib1CiBM2VnSIwdEjy0up5g1lru
eEqhGMwFlJgNE7EsN7UORmkbRDAcqie1ti11cNy9isLMZ5VLkyV4scj2PmHbRo+d
0g6OnYMM7LOyQQP5L4Lg85zWRvAUM1KLEPXTKaGUwx46fWdehAfXA4bjkIBcPfUf
5X+atFavbQ5Vh9gyBetEB9DNJvIysXCYeKPfKPsAJ7ZEe71Sr9iuh8nNuH439l8L
mq5Y1R/JeuAp3npuefvnWHv1OHK/B7+B/c80iyQHtwOP6GZ5/bQ98ZD9PW4LGIfi
wFciCkQ4tsaLyxfYUGfhMshGnBvu1OWSwFm/ds3fiLzPUABAUWvyk8lpDH7zJYZZ
7+xrqSkvTukI0fp+PmgD/SSUPLfIgE41mvoDiOFMD36weN/reuS9lEgoQ0Xo6aN/
jh2lyU3VtwEZT22EqZPhALpjlQrcS54QHS4AuwNnpnPMEV5K6hbxWOuIAgh4h7GA
X/osC/fSpU3R0j3Zh+k6x5l9/UI+x98B6wqLM2mBj2YBOKU6XvgoFGkaGcDmohgQ
51LTX/pIA4I9JS/JD/pHNJuvV6dSbUMQCDnlT1phvDIKW/lVR5L/QUqjajRoi68S
CU1hucg9Ml3okqIrDMBAwtCsR9kca22woDyhWZ5CPjA4gnTdAIQxFRwuFka5Z5fq
Aztej1xPLA71NO3dsSsBCzVaMwili3oyNovlq69Lz8hnJjdI9ilsSbgJ61of7rUV
9xP0h1ty/7HGDcD/Q7US3g5Bv/5s2wEGRjmLprCYdkUPP/hJhD/jh7K9yl6a9HuE
PzN5TcxB9bZusJdIIf09tEodlra4SVVmBTelcm4hzxfcLSfiI46Cn/ev4yoaNhJw
IESCFKzKrzAS9LgTE2rv7To0Xj+aEr0B9Axai6y5NjJICid4v9TaAOvaGrGCQrWZ
XUexZLQilDIkB39KVGXePU+hNdAXjgqERoovtIIVJC/+KOUre1H18AQhqujRUW9g
TyKjyBVoEd9ohbbyo2g1PQVDc76Cxh4xPYkRNO7ROOZhqdnyxysemRYgTfmC7pev
T3l14f+ilZsE33ah7TX+ITT2kMO+4yakDlRW2B+DRJwMjNwXUJTYd5byEqbyZTWf
8EQfB14ax50fiUwC3nvSxJK2jelx0PfiQLDaNcQsfLy8ZS+WWBZDx3CSfsso0xua
pJrRxMI7JTWoiTfB3RAbpXCe2vTDEZTb+EahWDCcIphAef4am3NFQ5YM9jsdRnUF
vgYRtOnhIE++nAMOykR+lTbkJUfnqMJJo4HSwVi3BmpnvZuGXlb3bNZrdH0DLLwA
XSQIpQoGtAncQUC0NV5AhNcw+VctI/yOudzwBfWMBDFcUVhR5vmUu+/8jC7gge68
Ra4wsYgKy04lw/DsF3RdaMYboHivYI5CRhsPseEr7ldTr9d7sKCCaawBG2Xc0Q3M
06UZj+tErgLKfbEWklWrhDOt09RhVcbyf7clUKB+GQomkd8qQvQGEfe3I2bQeM17
psPE5EcGxRtbY0lJ3spDNwxfrRF7WXqdN6BQ7fgnKrofh4uZ9iwC4dzteMmzCbdF
Vs7xFQ1AidyamQCwzFIXU5zk7ZTlWUpSoAQ8LJXi3n6hyuye9cnCkpI2mTbNOHIg
cMxyxQ2yqQI3vVRezcNjSxduvH09k5T2HJRyOJjL2nxsZs2vw9WspD9MFaC7lnZz
UKvpOgp0E4lDGWW8se5mV5n1nHubZkBr7XTEhtG5yQ23vHy+H+IXfWLMwbwvNncG
Ocvm1yRuXzVZaOMdnd7RKN3lrfkbiyA1zx2oJdqzaT4zm0qUh507y1UU+E1ws24S
GlWJeguLionNdPor3zxeYdkRhHZovZNg92Jhgxuvu3QHbH6gXVDjqICC3b27vsQv
JHFFRM9wcGFvaRNFeo6Q8NEs5wAL3tDu3CwX5ajDL/0hkU7TyE03ZrJsjpNLMfg5
zeWBTnkLW1Tu2ApWdfJ2D2DkuGtDXEeXt/TvKIKPTGw8c7NNqJZ9rCP6jKN0hxzz
sRCXhHH4uAQxEtqBqqVXgjoR21Z70WISKiNfxmDTGoVoP2ntQQnDJDVFhttzR1UT
cwcX1CBc7xTwdra7pIAAu8T5+yOms+MDu9snnKkSVugXgShI6Dsqp6aPKkuf17G2
Cf7xpJbynTGzc1ZwZGx0vcDD5KDVTNTwAieREpgH+mVnAtb0ueC9KyilJDKPRq8h
l0DdUQJMjDVzl/sC3IE88RJ4KYpb7kod8PDJr9o0oCN5KRCZdfoBJxQrx9JByLZb
2XtGmfqeIDW8Q/h6cKet08EqMtuvEQu0MmXxC4sDMSULXQ+QiNs2pBzWJwfoQWT4
Yw+LwDLQHsMgUsgxbG5rN3FL10kg0/SFmo/W959cRxX7sDh3eZ2VNmnF/7B3OatL
poE2BY9wi5oiyUcsSA10OMwlpws1kCy2C6XZuzs3PtyNzdgcWzDFcbF+G+BTqAdY
Jivzxg3JbB/KS1MVBwwp6XcSLRuxCzUDMBj0zt34E8nOLZuKNlPv0RQc/8vgp+kQ
GVc1UKuMNfoCgVd7E+RQr8xD390ghtaI9HJ9AYDkl/JklUXmNJf1UGMRqvz9h08U
DzqZdAVLpuUe9dNhR/INwxrEwGcdDbkN0OD6OPJsydjjNBj3Bhpd5o9ULaxsyKa8
fZZ63eheaBVjiWmPXXuJ3jQVRz336IIH7s6yLWg0e7Hj8bVmE/GnQqwt9q/MpzGx
0c/oVVjdvS946cTZkfWosaG4ILvtVfcTg+LePqmw1rvJfLTgN95O+rCQBHnzljpK
rnx4qNBAjwB9qFZNcaC8QXdLvd6gu0MO7o5sSmYMz2hK1B/EwRuTS/J2PG2V4kvX
YCT9vSBFn/Hm0UdHJVWRhYq0jq/Q4qJPRLL8IAqoeCf/qJ5e/UmgibklpSgFlJHX
isyZCk1FJYbyWnHhLrBRgJuGWMiiZwS3mEK/FqzN7029A4THW2jJQ0hLkipvSHJO
Agqqo/soY1T2K7xI4NEfIQQyeTynzXEHXZ3lm3aiUD+eIs4KKYCbWYcCBWhkB+ew
KwuHaUvEjxSp7M8WQwFkpg8XU/VxLrGhKP5bttVFBkPBF/odo6S42vtU3tkFYRlG
By4x137AyGwQnXbXrpaTThXepxOTKpUqkfRQcSDIizTvRNmoVSSC/Eb8uoTwrcOq
yf8nA+hBJTd3irk/8/q9YSuzkl/xKW/ZGNmtqkO3jK+jGy4u+Et59GV6TwVpK3TP
lRBaBMvR/D8HoHMYkMDn8hxlfHkg59Wi37jEDmVw8Qhxr23sla1HmCo3Q14baQPp
r/jZcsxMQAWR0rgEtNp9qSU4AmZmyTZZGgBMvjw8cFGmXwDQFJMbQZb+FDJbXGJd
ePvWD1yPoBMvOYzlqt+WMnw8i7K7duxIfkXyJwYGzdXLw3hhRHlT9bIpG4gvkp0s
Z/TpJHtez8nzh/J/iVKJ8ROHx0W8+S5N9h5WB9JtnvINyti1q83U/2HhEHbADmzN
qKr9GGDs2axL/x37vsZDuckljdXbRQ91S/yJYguzWoZC3DxNzpew20TbPxb14kaT
852E1McOM7ID1erb00ons92jJdmMSHTbXY/VPmXPXDPU1l7MrR4E5NSusa+JzjI1
dPRMkdhRMMvMrArCVEM5qae+Hlz1mMDsehaeKblQ/K9kgIiXLHWcCZahPLhLKpnk
5RHRRVsu5XdOh1XnSWmgxglkgHWtQq3wRRT6FYVMbC9KTh8I2aVck2bWSa8DPffo
s54l6TzKAQL/vTkje1q0m02Rf5UuwQNo9ibc1SzuP1jjGcJPgNiDI6U0ri58/WGj
lMA753ujrV5yf0fkZxA2DigmA/yPs22zxj1i7vVzwZ4MlKZIT0/0ovoYlClQn3l+
/37rHIOsan3SCQQXXTqa0/FQTBWU2H24ukYXWzgl+mq3YUwwpTWjhNriru8WZ6jj
3dvXYvqmXY6HyFoFZey6I9J46G2wOCNpL8JsIYBQhAgT4cMmAIhEXl03/8JjIQQT
wIXNHb0t5Yr7E0V8xqeb/d6730z8EmWVG33Uk/zUQX1pvprLnXNuwC724/HL8VG+
DyMYqzO57FtSDel5qkhZ4pBzMUgZkvNpAc3i2LtFdXSRQYb7GDHDYM+ZbNXSeLPk
+XXB/X+VtMMg66GBR1E4EC75NZsSEi5I0TrVsyToaeudWl9e/Kj0nBpqpgotO86u
p+ZKKF1WsS1KwN09devg5+pp3OEAhELaYE3DoDFntH+SN7qV5BPvhc2m+WXiv6Jo
/r0DcS5nzkDrwvJqWR8kPg7VwTQYt3En0PR23gCKcovOWXG/m13sqqJ7fRjvVhHk
N3WAcZmxsVTzqdKDb89kNvepoI0Qj80v+OvPYADFP6+Yjs9Kfj7ZWPsPZ1Fh6ECr
9Oq7vAkACdEr+sVXtVW1esC6jHYEuk+uGUzJi7QcdvHrR4ovdNBJePKn8rQuteVP
7wjhyhmmTDCouZtFyIvXJRZhp79x6IO/Qm7l/2rZf2Q/w6mOjnT3vmp47Otp2okp
kDbwwp3s53dwACsknIdedOVMj8okDIjcl2/fFi3HQIWICMAZMmwou41eRym0ozEQ
R9Pd/pf/WIM2BwSLas6riExOgPm+JiSxyWJR4/1EuMot7szIvbF9l56Tg2bBuSf3
UsAFkO8ccBDBFrCv6pZkwByamX30XZXjH+Yg1ie1ID36/fkWt6ARkcSbq1cin1Ru
A4CTXf90nMrqWW4zwfdfqbqUiXXH582EktSCAH2ck961NTL4GPadwfrP/o9Rts34
/2Ir1wFr+KlMbRfWBIXVodBzn0GMYRPOkYcdNfM3hWkSrr27bUkBhbZl6Of5PM/k
Dtn+xy2IuP2iP8762CDW3jTFPFZOUmIDdpYMTu8Pq1lONNvEgxLkEc4k10bSqM1S
PcHV37OVy+X+IywmSyfKJfo6XVgAnDZqdn2IvUnKK5LiNpS213hOugPgrGbDs2G1
Jyh9W787Kuw6TPrnF3ZqWslDqJLp5djLFz98BE2wDyWzPuHEUlb6iHgETdmu6Usz
JFSpZNuj60W4R77SI/EV3E9BJsF0JPNtQynilHyc8tpEzJybGDWLYfR0TIF30e53
koW6nzSuXkMMyhbWvPqjXP0o5y9KwnGxgQ8Xtz1rH/dQb5sz6/BQ2IrBU9C8VzSo
AX5fBQQ6iNSMX9gU1nNFq1ghsgtGkZqwJDf/dRVEDs5n2jnOcmStSOj6HysSEVph
8b9Z5Gs9yWJvb9IothYsNweppwowhRjal1vzWaEYfcPKD9WENqKjokEBteFcsgxV
XAuERiQ/1eC//KwNZVAlEIBurKHfFOUM3q5Rzvn+QNBM05sdc2rFsfnykgW6qwDq
NY1GQjutOIidgAgFJl23aWn1KbPvd3Oq3b//VF42HDAoH/uyRzNCANxITxPnKBAX
1JBlEo8Gm7zbxJEvI/bt9TogY1Od23yOJaL5UTt+ib8P2MD2z1EPkkgYfbcVb0d0
0y3zqPzWRaEi2ibUjMi92WR6MHygUghPxHJKza8KEvC1/hDYhMxNAbId8++Rv0N1
2kDYu/+DpJBcUgVifvLwHPflTw9kZR9/jQpsrhLTBD1sXjOZuwMb8lk/4k0oU87p
oemZ21dc79q7NK0Ao6A3XnDcd3Wobw/5lzaNna7B8u2N0Tmdlm9fxO97FrddI1qg
IVk3PYaT3Z5himGoyaFn7jw1SFW73Y3tKxVrjw9HL+qrmTMS10202jV4IelEBfAU
4iSB6p5DE7klK5TItZzVsr8GGgEUTlWQia22Gt9z3o5zVai/hAvezteprWqpi46u
uXMczAyPH0HK+J0xg1fKuJT1BzwdolSyrEMk837uPIyq9i+i/090iXP/QhKaThqc
VBYcSrNfIlJSZsxQAPkP9AA9EdCpejhBet1w3so59Vg+fN7ajehgeTX9+Dd2HlcH
79WsDESSvrV7XVpWUlQvQDk26XiwNfQ0/rpLmDZqCMjVSy9atEosWkHfMOtQXsJ6
3M9GWgUxGEYaGad1FARkPmmKeQWIO6aqExYcOk/T2i2/+OMQQN5YphOBBPsie3Y+
XbeBELAipLm1TwTD3ydT7DA+IANV84YOzwliVwo/m2L0JRkRnjoOdZrXlj6jtulw
4yk/eoekAFhV3DjVyCvzYp5ybp0zgvNaxY4zeQYC1K/QMXQZngeBJ9SZ//0iv8Mz
I/DFJZVZgI6bkSJV1xhRgioMj+uePsP00Jw9/vYuXcXYMeFIsYB3ti/bTbig9N1s
xDgwcTBbpROMxGhhXCBgl0zgHMmoI3NP5KxeaVuibb9IGGWoMigddqQzQ4EOk2gl
NL+B5dK9jTmsve0cAgqIjcRVjOpslO5t1axFJnh21+BJtbuBIVt2wx1JCst01oZr
fmK8JoMq0IZf/wcRcJol9SrXTGXiB0Ne8XldLFGcGmltB7Bjs5Un/GaaM3+MB5+d
YpGs7pqWH7FMeVLhwySE+0Z3zaR/Y3HlaoxIcUlJXiF5R/Fae2dAZf8fJoqpGPo7
sLBFpSpBvNuVMcG7e0ceMKr/8U81jleWXI99/C4AjoM7PKQ86q+HxCqes9By8i9M
7LbK5mUpt+pKmU/VhrJzFSqIKrpSwT5eDr3iztab0X5W6IBvhI+Aw89rq43rpX5Q
MKj+pOssr6IueKk6LbaHIveG0ZM92EdWfG1vJa+AUZDmFk2rrtz9KLIs/vu0sM+P
0CMKrb+BF5gwqvIGhvkNrrxU0NYlfgEsaE5LX8hCUjqWqjdlKep//9H1nEyAs0Y2
VtNs3DL57SkfgoiDgo4qRgLSN6F9zLxw+4vhADi/5bFw/LgIpgMpNhSIcAEIBtKo
BcCriKl2cDdZFpD3K44qFcageUBoyo4/871BD4J94cYvz+MmxLq5CvdFM12Yu7AP
ZU0sGCuH7jobuwa+Zmo4aLpbf1GaWTqM44ylvb3846tV5j1mFyUe4b0Pm05Q7ATd
ZcF4g5vNInYJseGClD0mHhijVTyfbWn1cptZ2rYlh6QYHlJb55/t9ORNhiNISsE+
ewzbixOxrD3eozTLRj4ZSbNzPrETbMqSw79Ep+EdWbAhHBC2dpsE0uJLCUnesmPr
Pk0O3jNC9O3pFRQ51UyTOmRYjqpzbs2+9+FtpyBH1ClxF3eJuLKpHXHqJGeedM37
uGjLfqNKxd5UGvUENtthyXJeSXOHlg5Tc8QCmBc4B3V2i0hu4GEg/CoalmVcVGS5
dM0itwKyo7TJPKYeF3f/aE0ajPmPs2su+rBdOmz0XD4ACZ1aztq3pMED5TkJYM44
HbDHA7vsq7WBzSgR7Abqj+ivIY2gh9FbTM0i+cUnVrhS6wTOU8ko6I0hkeOV56Dj
WA+T6gn6kS83dalxSHN+R5kdHcY9qZL5zGWc2RcRLbIsXye7UVsOi0I5PSROPRKm
rNtvRo/JJD5PECR8w3ea1e9vyHNg1hbW/TR8Mpb+wbNDvzESnxIDaFOSp1sg5OfP
LyevX3PiKdFfoW9K6S4YDLLpkWK96xUE/QMQgmz1n12ojBPTgSvVmx19u0xE4rrr
AV+v8RGe9u8waoMnM4ggbDXmXM+/l0UonyuwolCJ9bz6sE4nHzTdjMmjh4RF9DfX
dfudjffUzSQj1xW/d5ASa6CTjadvqc6TfK9PM3GK69RM+q8Uskd9O0ooLZIH/B5S
nap5UO+3EtjjpdVTW5mVivd8+63IBZyLHgYknb8VW3phS1dJ/HwhMcZrOTrVi+E2
pK7MCgWnFEyAb1xqOiR14ZuMAvbrheEmR2nAgBmb1p62AJ/VSEEYzTN1PQ7sN/o+
uS4NAjLJUUikZ6JdvXYZgeuVAd2UH+v4XFu1TDuc62htinfkY8W1NO6ql8RLgKmb
MxAKvYsy3KWcFlz62zHLApOYs7KV8WQ7Q7Xn8TXv59gpfagYgj27qEx+pUVsV/VT
tjrEh0//St4OGXGFYBf0Ox3IK5lg2UsjMqyCRf3u24ljLZ0EejWokjRBnfsB5Mjd
9ky74IcRmFE8Tg6SbgwORpPySbuN8MBzoOQz6gpynthYAECSgLhRBFgcNF8CuRv8
t7Y8emDj1i8Ni8+6ceEtMkDiqmic9/NoGBjiBiL4RVjANLzNdJR0XCcz/wEmcQn5
9iOTbPcFkohPm5XcvORuCTz4IL3XCWRvqr+VH6MlmLKkMY/ddpOrowiOy4M8Amiz
CZut2KHdeh4ILM9qEuDbDmyFKmnusNhcGS7UQhD7zr6TpqFcfpwBJaA1mqQnFyiU
uZNOP2oSd7mZ3kaPxsM1ZzJ9DFf0D4tocREEYZACVXYnm9UIDWn7G5gxYeE3vtlw
G0fmF9A+oK6fYhl/r55gHGE8nw8aUj9IENLgkOWe86Ar1iy+1ps0brSkPjjvQ/58
bfMXpNRa7dZWHBEcMcqvrj/QDtt6MQnGhWt+DuIxhpETA3Xv+6zBQXO/ARvC6NYf
YqVAVT2KJCqetgYq4/pof/SIlcPlIN6qMOz8EGcalbvY4s7Cu5QBbe1b4dtCV5jD
dABqKNVvxxA8ZXGUmd/8cr28HnCfimnuWUBnWJvZI3uWerbwd4wOcmCyfTPN+6MX
rMJ9G/zQaApHVtPdbycFrowimMiQzZztsRhrGDjD4ZgEyKBVMtjU3I0GeIXD5kXw
KbXZRmPewLrWaksMMDSQhahQBh81VKiU2aMLtVlSXW7fjgNbgFp/dliavqjhWtce
+zto0INa/ud021nXnFDym33Xig5TJ4xeOWiK/oR1o1DSOBFcBnw5SQbJuCntBtfE
xWTC2wpPbsnpWcaTOkv8a9hB/Pe1crmprg6Aqyj9iH00HCANShywbAPESiXinpYV
erM1t0lEfMX1enUpKXCxo58WP+4/O4Fyn/NthyXPUsopA9kekwk/bwiL/z3bf9A0
Gp0ms7FAw/JOxn3iT5fIEhocpEVK1WSXLtHi0Fh3hHyw/gHyWOpj2qiS89sQoxOQ
SWUSmOptoZpx782WMjHvitVfARPHG3A9/uKSq8fXBaRiBCgmYbZW7/ZUXtggi1sV
kge/x50UCvxsl9nHSEi6y1fjvn4lSFlRX3QfXcXlXOa4nwHVZEp8OinPNAjx53xY
XpT5xMHMALIBLe+us/Z2s9U6KBSW2y849nj0KbCisV3b2kFhRsIcvGYaMOtCoOSp
dhiWXCyw9VbLHRFFbezF1Y2onBuOXB8M2QG9YEQ64IyquVTliKKot71c1EzgL/Cn
q0513Mez3LiMPwADJeC8RIm7PMZ4AiOA+WC7kGrY8L+WKAMvN7p15foyd1+O5nV2
PKOuNzB8uLqBGWbSfwjDIau/dvt6jm1sPw9ttHSZ4q6GDtHbGsZLLFT3j7kEWffy
FcUpbNNAj0UP5Fz2LSp5XvTKr04zgpw46aBFVm0IeXB/exM0omR0sQ7ByV0Qcnwz
8lb+TGxHGYwr3Nux5ZuZ5EmkbckTBSePxUYGqUJ4PSRuWlt/PN+Bb8rOccQFfIxu
1HZB3fpIH2Qt7sDoiKMuxM8u0dxal1q0hNndqIYmxcvLfA0m+JKlX83OD9vlxzZh
XXuS1owd1YCSGsQuryOBnyfVj5qlv0p3zzLjg6mbhklq4+3MuVAOAFemRQH67hYd
42+IIzBSvJb5S2Stg9VB1c9OXa4RqsGtC/lAzc/Wi8zq6flRV8WZVjyyBvFqahA8
9BUNsBGD18+xd/lwQec6d/SPumvlpz2AOG5B4eJR8tWtPsG3pEe3BY4QYc7tOSxr
FZ6XGC8fYbYBNznpX4lf8EGadH1JffRwhnf40PODESr0074iYAlfCpdT3bnPAMMa
ElERaO+VFmYIytaomqbm3M0tUNrbxqZ6OX4P8LtJXwcjpELA183WlShVi378ZDuK
kjQSvnFRkqqXvDT+cZJhthw3dpwuCJs+WnHJ+J70QwoD50fLtjRzGYgUvXOzF6Dy
MtmL6eG0PNReu4IongbQ4ZFd8IdO5cDDIRDI990LFVSi+XEV4LrOo0SXfSjaofpp
s6AkcM4RYyoIOsBJ1+yiLqVfDculZpJ1jbiiZZE9ikeY9XEmVz0h/HQer63+LENG
1EidaUFsRfij8ruGC/YVv6oBz8YqeW+CLoAIUt9ghGAfno9AzOlU/CWFeKLXyAlZ
vOg3lhZKZmmIkgXbdynGyzSmbIWM7hiqOXX+7wr1m/13ZY2/rc1Ky5/xCF340ucc
r5nAg/XZd7SnMqyfe1BZuAQTPKyt9m7cgFGjVHholiyrXjiUcYriUitRjkT1LD0o
dLbal7ryLQ+X8Zcj45YSfzzRsnezpWblgkBTgEcNvQE6A4bF19ZV+qqmXJPdxFxe
PhVGv2Ho98VpCswdCtkpFyefTg9ETnJtHY2yGq+0/VKiu7zSevCHUXRct4UFU4tX
JT2IWMYFJCRTfs+03xkWGwT+oFtNYWydmgM89gl7zQfxkYBNt3rpRhuraOjcrnZ3
JYf2l9oQ3/7lmyfGd8mfZ9aDCiCyNruMRXFShYSrEot9U2SgbnxQoG2vCbHElLeE
EK0AzyAFmxZImPgzR4uB4dA7Vi70Oep9C3IauDtc7z2hcul0hhZ6nGJ+11MzndFM
DBzoYCprNt5UJ9R2+GDXFEcKLyNszegVy+Wc7Pl3bf1bqs4ek/ePL3t546POFluO
ELs5eRiLC5tkcJvXmH7L8atwgkLOysEWhKzTHnISbY1W4XMUU9zYbl8bC9/ah/nX
Gezlx+ZIA5/2Lr/c+pembRlqqINsvJZDNrSSRb0IlkNKoHRdLrrQH9sLw9jjz+2J
ZLjFy8zdJtgJXhaKxsZk2Qhe0IMnd5kpuhENAah3MIMjfANMeQhIG67ziAnUvTSU
ZxyTatrAt3rXZl5gZiZiVs51xDzIE9ngkCIP4jlbkIbL08V0FGxa/IyHDuolTnE2
ZgKC2QTz7FoUYeBcpNxtBxdWaqW8xKC6E/mJzQAIloKQlplz938H2dO5eGECEaG4
v5hKuWtlnldKyF5nE7GlC8BVzgwN5pCPL2ehDmodpr9O7fgNXydUJdUW9BDnYm47
TlXCM2kGBPZIYPFxvwW5bTs/n2jXV8bTAQ8g43DWMriORjHu2v4vf3PVzApyIgOx
s2IaHzlyPQNbhYpPXRvwkIdTde84rzVRzbV4S/AIYwV1WYE/53NmEJ+nwKFVvkRk
M8qvTk8FYjl0OH5Dpx0HDgC16IuGADdwwAKvvCmnd+2QMT342DFpY5vP08NtaciV
RJPy/OTo0d5vrOA04QmmsLbzSnRvx8SONRuAm6Xm5pZPZ1YwGMtCiPjUAiQayJ9E
bMObK1o28vfYIGX3X3wu03W+ukWuutYz52m4TpPuiykNd1I3CEgr3BeTNN3TGH8o
nTfcx1P1XqUqNt7x9yyGr2t/4KQPHqcaDVzV1VlAJWjIDpL/jvMOQtdGxr1lpI+u
uAjfEk/5mfxbxK/ad9zElSmMiLuQTdK5jtA1rF2UYToeGdmSnSmCdQrbHR514uAi
yYQdqWeO7A5KxEdv3D7BnOHribvF1AQW9Qx4lB1gIBg1IlrfwlwLMTGRxoAXLzfq
nu+TtAU0PyHtevysMSIiVbm4FQcz87dDZLkmg79ZgNzmK6JDynrWutnJLOeAk4T7
VIOkUAZjXKR5+r47RnR2oDWi347F6ZdmAzcw7IWQz9n/PweWfN2eXp9/0F19YFhf
XBZI8GFXQI0UlW5S14W+5CZjQoRdyIoDoPqRrleuJZR+7xEslPfiaTAZ3n8osutT
sV4bnjGsCWdUBUSwdsPbRsLNsQyYtWcoIx1nvUFpfZKIMeXRM+Enr9bi2dNNrexA
BRH52somNdF6p5h0USlAK+2wzksft2vFKBvQsF4hT//j0TUywrdwpzp2FG4NS01Z
Sp8jlf9TQBSkurYPNlDvGwQZ+DcK7VQuyj4jyEpTK1iCmOaD4SuvIhVPCzpAzsuE
7k8NgUKeAxMNhkaKErVjCavp/VOVjzm0TKDbaAT+yyKG26Z37XN8ayx1dcT9LfJC
AvK9kaWZp6c2wue3JMfGjNriLCR2H2SCYlDs4Pin82KKLrZK2lfDnyRkYjTQgzZ6
far+yjc5MKejy7efaXQz7zmH+oBfvG18FhD3cBYE8IWnh0bXjibxG9bIHD7WQxHE
x0pa3ToB5YKZlbimoV5QgTV74HzAqThuUqYCauDX9F3fLI/UU4C49/oKrAH+Ezjv
sqooyas1lCOugqg5Ju7j1vFmcIUR33x0cWRzfslgCGd0iRgFyPvXUfn4Qz3qVOn/
u6R+I6ZJ9aj8Gfd95Ad2ALJXKMRK00jCm38TwYOpkHSjSJvLfH13kSXK2n4fk9F/
E5Ob3JOAhEu03LG9pYnT2Ft2pjnTGcyDKEh8l1/cQ07YSGeJ6cpzIRx1fqcWpG2T
1ep1lx91IiUcq3ZXt6WhUNdUz/UETVk0R2YAOaXYDK3k6Jd6q21XqeQ2dpx819xW
7QbDCaJqNvxUw55gVzikUVFLq42jHoeufaWdG86byO14kZV0sV37lOYJlZL0YPVO
lu5tjXvbaW9F5X4nM/ajtGpXpUAU9pEN4Nc7C3zoWtrsg27kEhQAvoSjKSGRgQvE
YE6k/9aUw7h9jC3HT8EZ5JEM+L3KIiVc3Q+Loi4eDYskysyKaHCxntFmxSlOLbHA
NFkTzcQ5IuromUPQ/KtHPIAmWF1qGRnG+s5ZowG1RvD9/Y/20D+lTXF4qjN9tcNA
2gPaAuyAYLKbx+zMofTQfngFXhcUTFqRcHAKGFU5sErYP/OBc67udAmnQGdfw8DU
CaeSQ+7rhC6AxACmog5Z3i9354IdpwY7K/hpOWScK603nuZWEmYgeQc3H06lA0JI
n6XSWTobB2b47us4mHi8ve0t6pPq0Rl21wxwu/gm/WXAOQxU4tneykLDp2xaasze
9cqWKJ6nj6ERlQKA2XiEwBJhTgFRc7GXpwlt4NO2PYgwR8Qr2fNPxePUyvb4KRhD
SrDP/Ae/ZhRqWPCex244lGK2GtF8cAMxbCbPe6ntWXDHtbLqoTsfHZ0kN+7oyFvb
g/oeJ0Hft6vGdA96uVzH5mH8CSPko1OWmj8ezEufqsxnq4F3Uz3hCmta6jfqJ7OE
khdHUS0QDpZ6HDDb10PL2Sx33ZxHGYBF3E+gK6L8486uDh8cl28ALpmHn/zmR80h
KS0hNul/LfK3ICagz2yC4Um/YIx7OoscSLBXgLbY8nsp/zKkXsJW9Ey0Tj3cSHOt
Qkg/rijE3Nvg42wHRIZfa1QNWF8UlULFuX1wTdh7D9ilvIgwFvo754ry5cM1hTnX
wyfoEhNCHHpziOa520sxw1nxb0ShOFrDGCwWkNDtI8nXnIVgEHlAhXBWfV0OyxyB
iX64a2qpdIyW9QjCXhz5p2TadI+R1SoiwTasCLaW0aBmn58Q+N+VrKcaWdVolhvB
4l19l2LBS84y3Lys4YMXw5WoJvfg1NWgfVKAd8edEMEtydZ20AbiYjfEmUjUav6j
L5qIwDSyrhMikxtd7sbQwQefk17qN2h2t5zUhjgWzz14mdZB5pncNkYwp/uwvWgC
2vSkUZObdndnAVadlW35aFBLzhdOTUv+D0ObvH5YFGq+nH/NxUgnJoIfZnkfiy4+
tkJ7EWK7uGagu6J7kgbFtbdXJpeaGYAQgJq16t3COlCem+UA3lMcqiTmsmSvgLbk
8ldCvl7PrmaPv83OCeYl+zX2RvbXVaiG7/3xM2C1DgkUoaPeljwS3F0fzvap+YFk
S4pUqo1u2DGzATVLiHojdO8lJXzYetev0zk5MxVqn9nKHd6YDU+piyqb1DQNmp5H
hUAvi0ve0UhKRK718TthYa4L5uBgbEMLFnf2eUAkBZQsOd/b5iondEJ53CrTY7Cn
GWw+4a/kQV5mtPvZHmKiIwTQDR6Paw3xBu+koKmGZysI+JBqKOOppJ1m2yLIhjRZ
RA649t/pMcLqinC3m+6zalhqGIpDHJ5czu9cvcRDNJr4vGktN77CFhIecRgYWPVu
H+O1D4/8lkwcRaHTTlWEzImmiPSZVgNiet36EUtVi7Ln7TYjZS4NbneN8ImYBjqp
Z/3H6u1WG4tp6opxuiPuShidEpXkuOc1wBZn7NMZLP96eYyAczkQWRABm4gahnVY
uxxo2sdR6u3xvkq3PahE/TD3oV+WWkYKmoGoH3l1CfS8sszYrDF3Oyd7Qe07wrX9
Lw5P5HAiWwJl2lu9050vn1dnynIEIjK7G5GJkCusshYtuLiCgmBHT0rBihMTJ8Ll
4F7b0AHwPcoOwuN70xNW3oZRpbgHdh8Bmyv39QJ/yfNUNqsBkOHstb8uVZmUz75Z
XxBBPfk0RxZAEpLY2F5K63gfsj0ETapa9x7uCVWDgBW3AkNw3GX9ja/aCAspRFwm
DsLZ9WguMsbC41qcxCogYH9cist1mponeNvO7X+dU3CofjdXKwQHqaIabaNSwUDb
IqULS9ytWfwJ2bMiwGyae+Py/R1koDEp466HS+HUG07vCZYWxLE/0DNX4CVDifVc
Q5HP/NhkE8B5sGrwwtnuDYcxrTW2DKAc9Rg8mTCqRVhNbScgzejg+/r06jj3Gj7h
fOWDfk8CQHzOMYz79RLnV3hAad59a0wAxF6NjNk7nlg6aZ8BPwauH7qt633caj3r
93lZdVaCDYqxX6gcq4e6JMk+5+bn1GNM1GhN6F02EBJ3swSJkbZ2rzhB13BwfzYj
P0xuhO1ZOaWaJeSiw7OZEJ4JbC6hAZc2z2klYp16Rv6951Ty71N1vFiL1Wuq6UED
A7ac6JS26Okiy1VYPZf9CLZ7w1RB9Q9DsvQZy/w62WekxdxNadbgpqjr+n7gEeiP
qx7oiLmD8GsVkeBgRZbRE/qjAtKJMF29qhr2sSKQEywWQFYwE7J8J8h+zJ3tTxXJ
Mf1f5ZMaS5c59WpBuLFV4f+yhT5KXm4SzDtZFeOWkOKMae3PZoBQRtyb+pMtkaUg
J2FRPMK1MHIKevzDjYONzZaJh0A6B+HjTdHDIHhKI9cOeWyvDyz/aB4t+hYmkNHm
nSJjAKiSiSfs00g5IltXbIBFAXyx4XRWGEcdI17ZNVirO3D5+wke3cEm/XOvM57O
SuwKzB4VT1dd0NZJshZ9pz/YSU4J5WwzgwuBPBA999qpnMj8QChvred1GjXNeLfm
zFyHwLZ/YvvxRdlZbSg9R3+XkF29nskOR8YL7geFCSj3X54SdMhqbXlTtD9QL3Tr
IpU/s3xCPjq54l4YAEb3PXujKqQu/WFyVJ5g7lIa1DaCwOlvi2IsSMKjybR1Qa32
X8z5fGEzcdx+XTfTv2A60EsUHK75LagseoHqF4RgjrUb035lE3PItPhsJ+G6doW3
jHG1qSd3gI0Pyw6eMyE87csaCSnx4MqiKAeixywT0gkQzHu/0ezmjLJFr1mA5kTL
igvvAandNoA8LQptQL63fWi4sx8oDADF5/HlWJdyWjw6QUMHDz8Dlb/QE7Tg/vuf
POeQ0v4x8o0skI1FJjEQb9qierNf9M1Ss1uO9I/lzg2BR12gMx3r/YZvAnt62Q2y
CGxe0kJWvIDKZQyM1pGDnZ3QhBqJT2OAZkKJF5XdkfvoJf2n22CuPR70K8uxcqsA
gdQ+JyQs5EB1LQPUA0RPrVgAGEJYjMncQMz4oOhWkWxKyKGxl6kce0FJ5Jmcs2Gd
qNPlrfNtg4eOP32sJyVriEUgrbYyOxKq0MqNovuHQxD5ciZi+NXVCdonM6b8WHEi
icnJ9aue5LJJ4yicERftaoJAIVfNrS0kJfqV5DEXvEDeABN1dep7459XDqb6Y/Ff
aabZrNPepEGGB1OHTXov6Owh2J8p2T/76BMmGZLB1TzWj0bZ8d3/oIaYOJbFrEJk
RvMIPfkq0JaW3yfL/o0NxHalXa7WtoasajYrYjwjP3KcRf4bjPPMPRYNF9D8HQbr
IIzONF6xSKZiPrfIE4plfzIsYNAkK+X/AI048q1r8M4MylWEJ22DMc05xwtkcM3S
NI5PDBcqVdMAdYAMKzQRZkCxPDH3X2unJ39djGDKipK6Wze53tJKyKqDEnNpu3pS
j4wP+YQhTnwoq7unuGaVwMANnxno+iNHCjN/Pm8Ba2wAYsV73tO1MQUc5GGfvtS5
HmJr0/Fn9Eooa1dR+Q4xCwww/wpwp/D3WxwWUwalLIGPkPqKsQ+SOXf0W402fH/b
y7Z7F4SL8IR4ePB3RN3uU5O3cBwq0ycfVNfUoY/sDuyhd+wGZMTGhWFXFqbFhDbg
xiktftdtprkwErJBuzangn0ketalVh4M8QZNBQZWHWysE5v4bDe1nYntwAP6THEC
ikjAgUgTYJ/WTLVakOK1dSKd591AGCCpWZJkzTN4r9pMlVQp8BrO/YozS6hyyvo+
sn9r2WHqlDVU2K8LjUALgZx/1tIrhsiTGl7X6RoLK+gpIW6baCLTyOnD6e5ej6NM
On0AbM1rqXMQA97kPxm56B6WLd75tRc3EEDXgDWlgYTbAIJ4J47hL1hMqpLK1H0g
9Xol3G+D54AJGnOWWlanzOSzwt+bkzcIT0r6+pD9puU7kErNvpSvxnDVIyGKUIu6
h1uhdJc1uVPyXbjiPy1kOBRGtd0EMDvpA7/UhYvdw9X3DKMO+xjXnuARNgLXNuIJ
xV6HwojNgM7sXivRZUqa14pn5b9s0TbgTmPP/X1cwBBegh8itfOxsaq8rlDGiL5N
VJ/QDtflU9DQtl/kjBe4VD8GHUk+KZczAixyG0cTY71himV9vp/ejo0pupbeJmp6
tTVnfLzZob80hJZyUfeBjSSGKlh7YQsT3aNWhC1Y5dNp6J3NbApmVeOmL3aHYK22
v59S1gIf8AP+jeAi4yLzSH362w+eQruybIebs6Oya4UdBZ/8ls5h9jvtUURazTfA
l26vqpi+8+iP0+nnSpmntqlR9TC8eUv0GGDJIC7H7qOtXCYHjq/ZhTv/Q+AnORmZ
uJw40UX2PIr/vt28BvB2JX+pFgeOxD/P46rwtoBkw6dDXPeSUmYkJHdXYdzvfP/M
qQqe7xIEUywu6GzYPVgoK5gOju03Iszxcy1mps0Lca2He67s2jHTGwOksocDlJUM
JqxJjvzjDu8seqJEz5i7CE/gY09Grytk65CZKpR0LsedirEZJn2B55Pw41021Xfg
y9X53WVjrhi0RAVJDGGbkbtCbPGUtg1zhtQ6nWMQJwWYWwtADhkv9ahzdxQ9kXcG
YANns7yCOkexkGn/fxI+gYDoje5OprPfE0kOkqJhyQXDi0HQ7B9ql/8ocMmNlwP2
28E1uUTLl8cCm6RI06u0tI735yBb8RUfWK+xBxme/0IpWZAHhcZJzo/rqCN7dq5k
uhPgrjqGmHgMZdVAFR8xgBw7dIt0SHgEVCs1YdNWvPxB37xh+ncM5qc46MGTG6OW
r4K3LzTbwPBNSsuJ9myQ/I2vpLAZ1YYpW9csWPZ0hyecNfacGGke8gpMpxumaemT
6hJC5V/hfgkEck3I4Y2mDYcnJfPCiWaRSmu5KCqJVMrma7SSOBsS14vpVo/ZW3Yp
y43YBoRQv7vUneWzfgha0fYoaWbRDevpH0m7WhvUsAiLHm5MwheFlseTYOXq5Jgv
m5C10+W/tKXy8KMLZ0IICjIvfsT8A8ll6zfNfhrDyc4MIkugC+45jpZFzRsieelr
8LgzfV4vTZLHHd9RIGLjuxtM1c0RxoiTo7LylhTn2FnHgfArip2yg8Dvb/mRMpNk
eaMcSxp5L48XauceLKXW0lIM8RrMRyG5ZrLcvjovHvJfb/yKPw9jEy9/ntqCa1Cd
22IGNCdjFbHnEkckSg/6TyFQ3qG60YlDU0F+b0+oK7sLrkLENeEsbLdLjin5WXIB
j8uKDSifRGu/SxfpX3tex8MmgLuqaEEKULJdmsvAeQuTu6/ubckhPkULz1ntRTdp
l6Iw1WXVg9UJHn5gQ/fW8ehHyOt6GcWK2pMIJMz0sXQtVOAGmbavGwHZ9RCN5EAg
4sLAFETPZUzIpKgxF5Vpj4pHxujlmtdkZ7lqbEr+LtCspydGZmGUygWoU0VX1RbY
MSUl5hHumVCRN+H+gSRdRz23UnnEv5FhAzpT6JErEpi76/mJTgIQQxe52p2RaV/s
vvs1Bgg/VQfAI7RyEcVakJ4cJr08Sqz19uzv4CHYgo6OrUmtt9lLa63w1gNxX13z
AV4WZJAOyOCO6LYA8/a2Wuxh6JYk02HeN/zExoeQD35aze7pZRR3lodQK/QUO2JS
lqfIGBAoCzwqbgaardt+29Ubaasr49ekFOFvur/I9q7cee1i0DjncR005LU8Q1WC
0BZ6L2B47towRuC02RpiE1pBUDN/MlLn/SzjGg5Tf5fJLP0OJd/DTieqUxD9QpY8
NuYwcTlDAnFaWGjcumG8XG4YuZQkZmDrlZbbsZ0pqwTF74VJGB1nkeCsMONAiMSJ
jl+Zqs+55eEq6cVH4LgsAeAFD9E34FMbLhCzyXrYeqenbGiqKB0kydhV71cPLJIf
KFYO7zNybqjxE1M8o9RWZOvKKSsuHh7QWfhwV3zQIhNmKNvv3QZfQVH9ua79N03o
YDmQZCOsfkAWiCLLHUsT9QYBhLx24WJE+NfEkM6PFS69HgAxMUT3QjrwN2veaBEj
cSLP4uba9wInEVRzq7cIyFZwLBdIPvNT5LsKyEnTUbDVfoyi0rAT47SZU6R4Lcvi
87Ey1dfWNWt/a4f798BIiGdyGGztcbpg3EET52rrWX54AccyAdZsRfQgnkdzLRq/
POllFTusZ3VvHYW7omAFYGhYbpPE3AmbjALzIG6NV/7pRYm+nBV4aSF58MmFd2au
SHuAblNokdvLmAdrYLOIS7Gs80oeplC0BaqYRIQPtB28KYsZ8ztzXvr9AmX0sjZx
oOfSTOd6mJFSBCcaSKibQPhpGZ6+0NZdGXRrPkEhWBL5qC9v0Y85E0Vb3AiDSv5K
Y48gu6Wgw0CZA4XELVQZP5KmIjj00iNw1UQM6dW2scS4KczJedjwQnuzJwl2bz2W
UPIsYJLTUv3Ump4RJJAHKlnxdBE4hcTAd7cebrPyzX23WD3z+05auLP4x9i/rcP3
NUnBHIvJGTQlqR39onj3+nxaA7xDl3CCj3LMshdkxXSOuRLfLsqobxXFMQyVt6rC
eF3qjqUuvi+CNaMuEX+jpOCkZKWJN9bJg9zc2DshfCJiWf32PCH74sFpHULR1PY/
hdH9PuJJ5nmv1ZXaEKMyK1WP4QQtyeZU4yQGdTSJqcLrHJHWi4beY4IV/6T7Abdi
rWhbywxphucPw+ly0ByKzSdPFIos9PkdfBbF6jWLaCAjW7Y73rN/4kRuVhYAGwgr
OvF7O9pSfuXcJmkDEUPd36Ie2NuG01rWFbN55Nu4B1o5XIcZbCVOXpz/t4izcMlY
qVqjL48mGxBPduueVPSzGSy0SPqS7RHZA26JwVlLY95SX+9j8v9p9jWyimw03RYf
xtU3ESWp7yX416JxUpz6o1Zq7585i74/UUPW7SQ/1lbyyhHqXxMIylRAxx49C7xb
NJxWEo95DfrSXqW7psVEuH+vGmWdCh169YCdkJgtlshNyWSU3VsHzzHZO+A4vX/P
o/S6denpJ83Jkz27sljbR1m0mF3Hy0Bb0qz6Q0/snBlfZDeBQEZPPShN7IIkW74A
RUcMQ2NpG7Er1NJJSHCeiy11WIdlINnxTVKb/xY3b3z2pV9h/WqpcA9BTjGlmaN7
H63IR8rjvFGusJY9yHTkyJhxHXChjmZlrwrDPUhL9OuwJphxDGEa7OxJJcVeXTXt
B1RjfHQMGBWTvRMyAdL/EQHcsZ/kyBLNumStlHqqyIghf4wzIxQAxaHAj+4zn6eF
vc3/sDJ7wYQVSNA8b4Bw0tZnR1FZLBmk7fr0lHfBkLKAIhzR+iBlO5hs2BprUXuT
IRkjVWv5ni6QiW+4yI+03Owj9MKCe/ctjtQjojzppeVjKMFfEdMYDsWaMspQ3OfQ
8tQCHtHoCgyYnviqktzd3ozmfrY1jskwGIz/rAlfsUtJXPadNQy9hlfoJ/bd31xk
XjrWpuWcQcJiAFwsrBjP0a+Rq+x0BkguC/PhjLqxWOlNavx4re7lB9woJ8ClGi2C
sVdIKYz+/moaRHsTjajwCniBw3ae5qhbvGG6rfpMuwlLNgJ8Q+tf6AoiCFFr/+l6
wXT0MfnuNr3yefpjTzsEG8dDjkVI0uVU0WW1B1vlNJGNEHJAGwmxwQESTkyXTILO
E0Jbp4g+0WcIFOih01v43bLYP3uHiZ4sTIyEbExZy5/T6JhAWvgbZMTCkDoD0bsM
Mukne8MOB2MWMA2N8ZYe4wHTBNXQYFgHfNeH3Gq8JyhH1AnIzuPvjDYiul//tAb0
IKUXyfU6C9NrE458VOA0FNdTs1j44kT8vj4KmCSU0B4MyPIUpwte9hbcwVmUtYjt
Lr4CXoFMAOiAGMYW7Yh4/esKm50jN2mbu0B4/sxoDjVtuV9LTm53gW/cqcMQjU7t
migV5VSP90eOhqqaNZ/L1uEbKYog4TzSrI7ZH69iwQrZOMB5cvsc1X9K8t+f1C6W
KHYmZP5Bz854McsArW3USIiUtIjvUjDcA6PiGJuXScLJZjc4qh3ckKR9iWyqVLfR
+rn40DzcGPo6DQgv+7l0Lzrboyiw8dattIo1ZiHZ3DkiGFW2V3r+DITc48wrKKFQ
Zhg7eNZuDcf2TuLQ4jJcBgHvdylzNhRhDSCmOX++ZlPXsYlj/IkusatY32w3aiY6
8AvAauNsUkHk5oaa65t96xjMwGado0/OD43blbHQL9/p4uGXs2rPqVjs0oUDFtfZ
zjFUWFooSG9RDliN/HYtIMqKvKXb7faf0ctPus4aDaHmkoX0QYEO+a/i/Wy64Z4B
ZYixbkGT2b5b+wyWzsWiJ1MCzKJrxisgZNr55oLmTQuKxgvyR87z98cz+G1aASGK
KPQO7ComNmRDI3CykbhLwKl9iqLFuG3+AVeDgJ1NgkzrTZjxzOrH5D9XvIOuuWrL
CYaM3P3EX8CKDelNimpE/hLYj0zKKmoVnDystoO84EV6oKVTwVZANQKAFlxy5lRa
NOqiqcqRmNxeq0vEUKsmSVeWjigYBZ+HYYaJ+fKB72hjho5jbFd1MiOO8v0lLTXl
l2GcKz6T4a+8WREkWVcPh5XFkoVLwuRqhwTEysyaeTVYdrg6CtvOoVgQOVNAaSs3
x4C3hAk2Q2elWFN4FVUEv4Jrug68O5rF/gMsBbHLqaTFCWAre9di/v6sRZWxSvsX
R29qAKiJQ6C8OKtcvjAkVcNjBv8VQCPXB+UFoDibis30aCFulBfEKYdxdhq0CAKQ
Ru7YL0O9x6hDnTX1ytOmCjboYash7+CWLVLHWPrXqxBJM3ITq6VhAy0NseW7AMfi
qEeiDy4KVb+U5vHgKNXkPfLDXQhrFU3AQaoLoY6e4PNtL7/yb+tsRx1o9tSHKU19
3Zeiyf7JgSkSNyBoB4iDQTbf3kRcchuaYFSDAakQMv9WBwCruFgYTDN+Ykw9OkYV
wlbIHQkJHP7W3SwsX1hM6n1/V3D3HWTHKyxocIKBnFv5U2xnlTVXyaH3l/YnkOSn
5BKTnsnl5/wrVeE/0FWtoabfbmPZR46Kx//NGcwkBPvus9b2zgq6CCVR8YFBqtdg
1+qOnEGW/kDm2GZyEneShiPzhr9yWNx5ftzlPSa4EzrQkkwPDOK15KUO2Yiio5Sc
gJFmHD0Iev6vYtTsVQDh1ewJ+eDzzk1sjFXscTLO7FYgqwBZYuK2BNNnwAWcTNmU
ujm9EMn6xRYJkJk/wLpSHUwOn2h2MSeOXN2sAG6GlQtzZABqwcxcYz1O3ZKvGNp3
VtqvjGhEDk44g4lN8CYgflEmTHHd/Y5vZlqvZMy9VYMzBQ0bIRnoAboECTR+bQkF
/T3X5BBahDYWHG5gMSl+5/zTQtzuflw4cuq/tZGAJTNGOJHEDm4Q+o8UwN+mnSBp
VXezhsxfCoME7H1J2sHak/6xGj5Ipf4Ef7tl5kU8g7qfLsx4Xsnm6eLktjzCFcPb
KJHLJxdLfNItqLuSl9rI5m95Kk2bMThC9K3cmiMufqhNaWkyM8aLvfBwDx0mKCKr
MZrthCqrHWXJAfGMJ/Rehgh5xpKmU8oi/zrUNAQe4CYJ+iU0cH7asbSeUp+B0V2K
ClVZIfdI5VppcV/Aofq6DOpgC04FxFNLfdJtZYZVNDP9e+oXEteaNhne4YLPltSD
MrgrSa+b7J9Q/I8rMpni7HlyZnQEWqM9oUZm6PkpPi2YTZU7hkS68EwxxBF6p9Dh
c9x7UEr6pDkJxq0v6znHdeoQtvpTsgO3WIrYkXTatPllfXT9r88yhkC7W28WXA85
2EOcsBF4BiqvtXxIyVO1J9ZOe9hcWKVV1kh4MMWPVXFaxpCz24hNfN3rggFKbmot
MRBEzv2ZXF8nis5TF14U1Gw7QcRKgCyo43QnqJNpgLqoPwBiAtfr9Nw14YyjBbS3
iZ4ZJkOarWTnaz0t1xGpCw==
`pragma protect end_protected

`endif // `ifndef _VF_ADDR_RAND_SV_


