//----------------------------------------------------------------------
/**
 * @file vpr_void.sv
 * @brief Defines Void abstract class.
 */
/*
 * Copyright (C) 2007-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VPR_VOID_SV_
`define _VPR_VOID_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
VD8KoeuP7j5T73ATKZAjZai0b3D7AFUi84reKBvn3j7KWeRuMRobDl6S5r56pXWl
2cNh7L8npS7/xPYSUQOQOn8Q89M/XrJbb7V+FaTYn/W0lqiaETqwrIiNetiM3IAD
zy5Ci+8eMvelrAfzDUob7PVNppGRxdTrZJtLnNyZzj6kjd2tF+/bEg6UWN8AzOZU
0KAU/0zKjTTX9lOsF6e7hFY7lBLatsYlFtVc/CBOcCaGi862jr113d29/PE7g72U
uqAOn+N/XEIsg8vodb29WnzY3dWJ67NVgvfI7PBYB3aIPCAkU46oqTMZD3sXwIw+
l9Pa06INv17u9Kv4cZuSuQ==
`pragma protect data_block
N8eYS48sX94AqpesQSQEJMUftAKe833rVvYIiBs4vAbQxvwjBYCEaUkgmdm9hA57
QkHB4tVyLIQiIAU+yo4ReSHYrh/br+peZ8t272uRU7lbnwpcKXpqQ1KEkOSHsh9/
zYWaLzx4YUUMKeuxsn4MGBuIqv0Z7dfztS/XGep5oxBp4tnZkY1tXu/8T0m++jPM
JS+P7LEIRg654t6j3J79VrikiWGrfL4a1xDJgrAK3XGxm30VqXCrdFLiwVIjdMvf
Rn4P3c3AufAbbDRiNgzsFciys3GiXCAEkCuu8ngwC0l0NuZM6CglA8+s+uH/CE/q
r27Qyb5SMFZXS5UmW/rptQ==
`pragma protect end_protected

`endif // `ifndef _VPR_VOID_SV_


