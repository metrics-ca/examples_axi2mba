//----------------------------------------------------------------------
/**
 * @file vf_mba_xact.sv
 * @brief Defines VF MBA transaction class.
 */
/*
 * Copyright (C) 2009-2016 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_MBA_XACT_SV_
`define _VF_MBA_XACT_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
Qvia6MDnqygQGSq+h47pYgqWiIWu5EVeDPamwAUWFlrp15x1vaqbVwRN6cdxPkZ9
2/7jZD/nB1V/mQbkYYcU2NB6gz/9GOtMMQP1+IQr7hNIBclfr1TmDODBaPE9DElB
gZ4rqJi4AlbDfEn0sOZ7FS71Fd00TXjdUzkfG9Jy8D9e6JfvNlokoTc/N9Q1GZbh
RLN9dwHlxGAHBVVxfgGXJD3RviN4Y544K55GkK86LnHrihPCXW3xfuHYA/O4VRrI
zP0qD+2tdBwpziO6oPJMF3d9hFfkKUqtzf/SmWcs9HMfjn2rp4MZ+OyOylT6W96Z
LP9xepPmDu+AddvBuqxsXg==
`pragma protect data_block
m6YEeqSUiQPidVpnA9Dqx+tWwiwv5Awc/K/eA58PDUXdU62SB3/4wWgolQQsSPha
QCJLKMO/8kdvQWqgCSzJtTZMDtrnf3BpFs9TMDYzrlhSEcxuq1PjDv+6BYr/8//U
e24nFVFOQv18FNg4eDpufgfKXNRPIu4Weo2NK7SSSWBwxQG2Y9LzH5NzNEZoBJ9P
LaHXXIiO2F8tvoN0cPkdJs7JO3tIfWfOXFEj3u/5clehSPHU7xZ0E0P4pZirG+oW
zao0cOVy3VFFSKareNns3nDWZxaqVRmhkZYy4fs2yher6kaBdx2JPX1JtkoEcJhn
bUJHfjAk48FeVirCxQefT0cDRzsDmxwv2i6zioMimOG2Io+tu86T69HqS8CyCJeP
Xdt49p7Gkn05SKJf6hzowcBq2S15fcSvgPEZkwl0E6/+zkGkg/EZSYwLA0iwG+2Q
8UEUpGc8WZeWuVsiEh2c+zYzFdQfs96f1isT6KWUbC1MMY1X9NilSmtqb1PvoxSE
lhcGdXT3rDlqwryZt2PTr0zXhHrHJ8GFKowXqo2QVdO1iohfi67FEApRnwiv0TRC
Fvb6jXHPb0prqpxhSX9Dk2Ywq7gNT25Exm2JP9HQxiISTvxgJjRm0/xS7dwaujF2
TvaZSWbHmAY3e3i02VzjCkAJd74KE6NjyIKOuWOBT4GeFZrBiciKWZR47HeITNrt
QclDI812u7FOlkpYl2FXBNOuzo/ImKCOrbGs3vx7+m9RYzH+sHfKcTakSui2W+xW
6CJyciW+pnfH9ZY9cItw6t0AF8jqvXjqTMjcfb4+53+cKzDp4SmhxfOq4ONEtULc
mStovdU+a95aQCBtVLWh/YP2bGvjm0gOzxF6vEWQmy3yS9dRp++bEoZiBDQ8qDm/
QyQtzWFg4LmsShB/xRVFu4j4VSnpxLvMEJk1u2prKaX8Li4MjvphfCmlTOh0mqmu
aaiSfVc2q12xtV90PmxxZM0BTkFjlgQDbWHY116Ebf9xOLxixmr7uPUbug0UXegi
bWl2AxUSstPBUKy2LSACCAZLZVFekypE8wR78G2fOlJW9j28/0Zw2ksodnk+E6MO
Cu9GomXK/hoKNRKNFYbB0BWa9uEm7Hkl5ybD3k0nvPo7dtGWTLUvemy5XqEfBdYo
cUMdnl2EUmUHzZwSR+R973MD5ppYhpCFKG0lVfGC4MnW2Zf3oUHpuhIuYTCH6kx/
1A9mPwOsybNnozNzO4CIO+RuFNZSx38myxC1e35YdhhDwSRdd04Upzy7tsRUmr45
Ftmxq5sWVpdmPaERm7YKWD4XuHQotUv/SrZnfkGXe19aguxIC1O6bo7gLDCMemtq
/b8nyTFXWt6kVCcpYsTmc5qLfDr3v8gCUwO6MkLRqPmvGplUreWUx9cfzcpuUK/O
EEoj26AymvKfRVYQYqdQMgzQ4LzVr9obWEYlN1dq6k/PmwLnQ4FF5AzJSekHs8P0
3ec/5+ykG0Yog/HkFkQDaI2eVBm2xpN+RpbfxkKx/ESShApws8cKXyC+1EXSY+Tq
nn3ZvE2mgALoPp2X/SWQzoC1UQx1Igmc1ByDipmvtOKqe5hjgETlpkY7YXHbUGxh
2ooPiyCy5V+tNYBjMwn3Lk4ZTujFVWj0bPzbCAx/glHmcPDnr+rzy9uP1vOUntFr
crbZwAA85GTIAGEOQxEz4rhXAtOO94/6b2wYUdPEk2Ab9IX5FbkkDkLZ9frkpHpc
Uk/uNvcpacpUHJtnaS+EaE9d2Wqyi5J66U4m8X8O6z8vm1hpghXnPnxJ6c5JbsB5
7Dag5kZT5nED97J/ON3piHr8lBgtkNQAYHDQqPl/i6zGJT+nPmTmxIiidJOim/ei
yXR+cEtZ3aSpZsyVh0STtOD8UWnX8kHwqysRmuHXa5Bd/PkyM/b9AbkqJMIp++dS
v96+vtHQXZxQlJ+a/oIYnyfIMLHJmqUu4Sq7Wnjv/3+hpAcK6T/VG+PDTFQwR/dh
c9VQwOHGVegRzeD0SBunNU6qcpF3iC6ABEe7p6lc/Bo3w3MHdyy/CIrIFn/O9z3n
X2C7wvCLYNRwBbqDXoxaZDxyRWg1lCo0RjrzhLQktbjrmvdz9G8GhC/Zd5guCBwE
o3i+xxxjVAigNb0MtHi0fVv6KDKB+nKz9qYxq5SnEzlhjHH8ENBcwqO6YqNV2zE0
vDR+FdoFDFQGEvD+aFmJCRu/MlcQxA5hWWp5KtH8wDlyzkfdoZ4z3hhpaJN+Tt5C
wJaGxy8TKkZscKgimktU7SNYFCMXISq+2jvsUIcli2uUp3J+i/WI+fu9H0Y7gfp4
Ho5p6P0uMXG0STeQVzyc4pfLA1YuOkumBOFVOL5twtB8yUvUut/MKL9OA0S6QBEx
hWlfI6MtmAN6fjvNrcbhJf2Sy0od+kWWKQqEj/NqXsuLoo37v6Zc+Tv/s94kCvUq
paObc0vg34xonvBmXT2pPYxQhKnD41h/4R6cuVRbJoEAbvGjHIUTkTwMb3tO3nxD
5Bmg5uYPZfM3GVKPy/jJ7ivjn9uceqrfEQhOk1sGfBPp8VI09tL+KJfVS/uYvPlC
c37A2hqJPaFkl4sGXe4IImpc32yF5KErteS2zPxpCO52uFYR77ylSWC+VNWlnLBa
vJL5DlvK4+Gz4gh7pLl0C9bvYrRhaEvsnI1VyfTR2PGJRkeutcGY90xbhIwQGXQg
hThWOshn0qgMOBtkY0iOfMAvoiP/WFZXRfj+ClSzg6J6TCBHn2Tnt0u2zmfHmXpn
oZ7J2JbKA+SEwnUw3ZkEipfq65FSMlPzzXdeTndLNXrBDJsT2kL/rdtgjpW7njQ3
3y4nDzMnBNgG45TxlYuOE38WCgC0JmmN3voImranqV9QBvV8EGM9g4+yqAytxz9q
EBhTizJJ1BWvqXSxTkQO/2IKdK9I2+e18VadpGZXu6kHS5keF6h9noqmZgNlvJP+
7hgrsqE1ZlKRCYRt8RwI0gUDv98V1eME02YWEGHtfiQZVWKEZr/wRh8ywArjZt93
6ufhH3hn3HDhYCm0IUFMmyOBUVhmF1ke2lsMtO3QdonCecytzT0MvwCxuDUQT5Vh
JT1XfaTNCPBsrrZJwGRbruPLiU2DM9oYYxpRNz5UQp7/SNvpj4fO+J12Ax7pCKZL
jgvc7YxS0Z02LQuhqMkkciPanyG7gqQtsc1F3YaouO7m1aTxdU9kHff9PubvmwYd
ld3SyY/O3MtsYFC6B9XNY8n8FAf3hI4MjufXlN/qSxqIv7VOkoT37s0P0A6XFELi
ze645uhGs+npWgqtUWlI2gWOxuzWYhFV+471BGBhJVF1K3iu+kzYeLlVPYlvHrJE
yXianIYfhtWMyPlgLLUH5W5GkVlLjz4n+Sm7vg8JvaTToBRl8mQaLfaJUFJrTbEH
V4waqXKqLFQTei5ouJtKZBum1SmdaPIKIu8RdQStMpqDQfwD9MNY1MLjUv3lfyKZ
kZocGsg2u+6i4wMBkV3g5cqeOdgszMVQRY7zaKVPFn47mdQcDuKPkVtixcaZybaD
Uplb0TbY4z8X2B4QeyzxNFu/VJa3c1eZgUROpxzFqJJsv940AttYiDBGfHHK84zr
QrA5svdMbdAjAxCfxCufjS6O8c5ILEK8q7BveP4dqJJOCfJ8HAB0o4U8a7ZpCZh8
Bq/LKS1w2Md/2rbF7XDnx5l1kiIVGFVEsHp7fPb1HNwLHw9o0oUd7BsdDVW4SCHn
BbdhRByzp/ZuU5fGQbWWEobOuBM9zJ8GlyGKO+hUoZZGN7a5kCPp47C5Za/siGB+
RW0K8tYtGH9K8iJchxDPUT4gvY+x3BqR1Tvtm+IFyt6jMzf5nEQ56cXKDQDG59y3
L/pkihqI3T53WdM5aJB5sU/BFRSQllb/F61GYijEMJXG5QiHLNPpW53IAPrEQ/HO
9TODCPIEh9AlBcsx7nzC8W47U+YDxPrb8/TVeP+zzCTsNDIQVk8WF4uyA9kXRMJY
EbPmaidUupUIh20Ac0T8XgrO1E1+ND8KbyKwIzb4OjBkGyVhvW+UaoTLlz1mu1Kf
16Dl2X9R8v6QEi+pPSfJT5dOSbVC+3vXuXBidhGPzlaMdCJWWZfr8bKzCRCAEYiJ
qlEzoXssTWy9+JF1tGVHJ0HhnNWzUCxKkXMrizgRF+2mFPxqQNZzmWZ35fvZjV/p
cePUPCMJ2EDZ7nodATqwUQKuFQJgcR+XKBQCrDFrwqo0CU5E/zGPPJ6Qj6ishA3U
l1vnizRYwf2qwjtxOT/tk0l+XnsFZbxwroqApTBl69wigpkjjNgwgPvecWl9nIUc
7HDyi/SIlcbCorhDsRvo4LE1cWkVIXu++RrCQLj9H69gvCPEsq4a8DxvV+7AMNPn
fqEIUrdTmT8GdPL+jBSEZi7LLGOiL3oP0kvpic+P7qHQnNFt7to2nn06YFr92U+6
T2QoOVMzil5vGyg04Vhg3yfT/Ruks/cZrdrDGJ0WbPFKACynDsI3GkFbEgjOPEyf
H6jSaZapDrIWuMNFKPNbmIF9jZzQu1VUC+a+Rvyy6Vy/6xgw8SizUCRpJgqrQdAn
j9hmoMpjGUYA4BXvhGQL9vLv/GlW88WkBFwX0sgXRbrVO+YSWXDdQpDdjzGUYOQ6
4+Ycp8IzcJyq32TWNjdGhZHErp+qs0FQvs1YEKC+h7gHSySfJxa8szkMSMYQK2tI
3LspOrVI1hzn4nduSCsNziG+OB1PjGWtHNM2DMn9shObNmDXEwNbQgp0nYgMKiMd
u9qro2mFQp7b8SqtRU1FdwtH0O+reMEpoiaYb/kFktryBHQA3p/S2ei991Gp/VH6
ieCl5gKzj5+cF7vPHHaGEGQ3HgXrCAfwYW8+waQ50srwiYSELmjft2MhjdIYImx/
FD1ShhU+QkUPTz6QD00vCPeuItHMR3E53W9F95pWxcKXQKEJh6PY159VfUxzMn6p
ju1KaQfui+fgh2YQ0GkjnSNLSsyI31Mh90w43RbcN87HRIhAAN2hNq44aOavqhHr
bGO1cNSRINGkwmt692dJOb3ljGdWzMOwYOBthOcmMbVPsu6Jqee+FxAlyiJdU4yF
7mNNuC4AGOVuCPKrlfapzl6pNLvZwmqa786yME28rrf7HxnPHQ0FrNa8ky0W1F+3
vvGp+B0FWXAVvHeenUFzWVRCAeHmnKXWW/vSokL8VcxrVCNBxCBEr8OGeI5/b0Dp
iT6Chi1HAPcBnmF5SQI5xfkXsioWA3XFOLa07qn7ufXQd12oRn90luAI4yJScvhd
YfZfUtCoTdyD7ku/SOKDLgHoc5PqJzA91SD9Ka3BcfI/qHvJbC1OOsXkKV18I+K+
M+DmVWceRGtUJZwgJicErZClaGg/k13zNTSsVKqEA/cTCScqUQrjqHsoK/4npZp0
G3fKytYjRzkr3zqtnc1WamNSTFy4n3jiKW+DmqwxkN88JVLe8T6YbjnzS0q5FaHb
cJekxKz3na6rG+luOz9t6IVWLVtPzXVdETbPy7H89JCco8Ayrpx5veFB/ZNG4ZYj
mrk01bTMRGK7n3yC1EtFOG12g2+k3OB97OakQzvcTKV8YU2EChkIxz6evYFYvbTz
dreaZpFybeZv7iQNqfJMxqMpEcfCGBoDYTSEA5rIpQ4Udins1GVWRKcX6g4BXpBR
+s2CeWXfvViRYbQEPVTd1/OPVoqmYpxVCty7hcBfxPCkf7semCYUbmRwwbPj8tSC
Us2p/QP0snNk6PoDRGOWpjb4lk5dPTzA+vDIYEIE8SqKITdQOjwHJjgyQ+p29hiP
fHewJqbFACkmKuTWUFTC9jvekd9FnSrN1xVfw9tJff0HXHmEBdvBIICyZglf5XeI
SePbddbMtJlHl14QajNx9c32g2glRE8WcQGviDhN6y7CyfvTJ9ntZb5nf1qIweQz
6bIvvHRgXYYXQRfOrXvfN49YtdNXOh0oZOV+Dz+2iiNu9s9g8Aw2IGj8HK3WtCJA
JHrriRzoV8kwZEMXzr06PDtPbGCZvOHGwJCtrzKL1RTBySG3F5sv36I0H3PMmlAG
fPUPHyNp/X+MLm8G5wRk4tuzQqwxoAMOfiEmFFulqTRik6Zo4pxRqmKeRNe4tI3I
egvGHSsAs4wsGVuI0UJpSDmK8jLC9du3Adc2jByzwZ9CHDY8Wukq2LK9tmY7AZmY
RMD7gYDtk0CHKSUwfQyf1NpQ8JxaB+s3Ezna+kO6eCfkedlqXOL7DBF9OZ0iBayF
8YafdQkaRVyhP4oHt8IIBsRWfqWvmTkk9Ttpmrh0S2hW4y0ludmrn0raltgPPK0W
oAqtDn4m6R1yTWgyUZ8pxWj4pw1soztPs/EFPHsAiwTA0iZA6+yqRPA95OZhmvPB
tax5yG13C+c2PHrtSfjwEFF2/NyEbQcU0kaSd5g+7jtuQrdkLofFntRiq49SjKp4
uJhoMOcF4seNkf3IRzowu9TUK5KCWV4QK/X+IA3gNbNuPnCwiMPDERRC0mGhxUD9
+5fAInNz8sm0+Voq40QsujoqER3oIuf29RqLgJPnoIu9L2s2tRXksx8vVa/kBvYA
fADp0SnBEOpySKSEUN6oDLM8GsNdf2hNr01eVuhA8XMk71JbOzh5ZBV40DwjKYqT
1n2htALi1XV1b2M/e9VUUhN4Cu4w5a2bQsJLb6AGC1v0OYf+M7ByActNc4dQ895y
GkAMsbM2rcbKjszAoy8iQwDrlJZ2tVc3kr5yjVkna1J3QXs4ham2oGTQUoeAE2TE
8akWQut8ixYQcsGoUwAa4WiEVKVrfBiX9pIBMNpQKvZwA06litFapbRwnfMu1hID
R2YOSFiTmGmXY3pHuLTzhAIk/dbGxtodedvsbhqaquhx742c5dDFMNAB2cD9m8YE
AqOnet+PaXMEEYYwUhKC8F6gJNVDWLVa4/TQZA9cq1qeKub4XIIMlG2gECrnWrrg
bb4Cz7v8gH01Ye5PkoFWaXFwdrar0IvOFrCryCubGgRVYRf1sFuqKl/7yRt+c8Ss
PxzC/dnv8y8SA1QvMweN3eevEAEO2MNdAZ7pup7ysXTGoF6z4SyyQk2G5uFS5YfP
D+0irtcW2EhjIPnf8+ruvUFQ814ThR31nGmmrOjRNkut6FQbFjcOmZdmvyF49yJE
N4VJiIp8OPKd3zc7fmvvfc51PN2WlZYulQOI+rTdr5BzC8vXYyIjALOgWd0VqJxH
VQp4rZhjDMaKJU5qGpuiAvWhtHwt0rhSsCXcTbk6rK1C4QIYoIyivUCEDMFuLkrZ
VHBWfp0Wlo2LZQYiuEPSOj07ciZYSAViUQyeBn9BVVtKTjwQfsBD0OUbttv6XNPI
aizWBQiEhRaq0IfKPKCdBPeUhXrU7DsiuyQYBJI0DOysjkVw7EOOGUeLc3/yVLbd
lYaEk1kSV+uog1T1RIZNHLvtSygzRdxfUiuT36vf+tVuhN3RpYMwmuyTFaaDNPP/
pcXZnaUpiA4cgYyXJtFNahr/8Yf55TyjDYsvGE4FoP8NnNWL4QFuhdD+1j8TXX+6
vUP/lt2GKPxIB+ZWONqZoYiLR+5/9axmsiJK6FkzLsGh4Ej9XWOj/s/wZCsYJBZH
SqgAH7xCiSgdj3DUcQkQ4uJhey4VmT/7jehqOSo2ppdytLEggxPno7x25btm1RyU
gCjOLo2I9k3ylIaCkzsdvwERq5wfW5YTFHU6BVL6UFXe+o4qcm+noS7IEyyXzckQ
cCemsl9hugoOKlkdbGriGZGoDfmFUqURaOTXvKTmDvanTQJv+NNMsXDWWexEwi3u
aPLJu45+5UgMA/23IZzsXMAh637FoBSxcH5LHd+bVD6yjYHygNpTLlL992yPxRaH
/qSeN3faXzKTaCLWPFQbbEfDrLXoc5pvpPoKfwnvaG8USGOhHHxPabXdIAyfy607
BPGqnYHhpK8WB/pQdRjoOJnbcBtISDQkX76mIoW2aIJImvuJNYVJ4XkOOivhKgjc
07X4iCeEwjZK5Ul+F0ee+jJnbo850UMq024tHPKsTDBOqo4CFPpOXybSwz93qgfj
l+KCqsc2WEvGSHgHmOgKO6wORdqlCauImoPiU7hx9gP7ufndzLuf0Qw4rFCTKo8n
X8Qzdg2h+NB3YBZa9tYa9irorUOrJPM8WiTUe62hCwOZeUf4BsSInkp2soev5Mbz
l9yidENMu1r9f4wGwLx7rG7CxuvxPL06VOVG5WymvPwAv9KVq+PtfYnMbJJXYRBj
P6m7y2Opcs3A2D0ngMdgFmqpm3gMsK65PpQKJwnBgkmoloq2m9LYYWOqwYjBqvsk
OYlyQEzY0qBqzZmHfiYat7yaNSapKUBUJXYkZG5ZG3HZfkZQR5oqcBgJvnAxWTjt
y3l0ATzwhZz/tg5Ey6rQRUNGsXYMqT22m152Rv9nu2JuwTWVJf24wLjrCUiwwX+0
dJvgbZiGrCKgUir0uMGg8I5B0eI4fpBLVrTGA8RpYy0FjPNT+OMtMWQWWoDgFgB9
3QFSlbu4fFcTA0PpNtms/zlNZ9v/AbEIrxe5g+CBPkrX/rPR3nIcopz7Qy3yA22f
6LSqb3MQjpIyf+IWNdh+aWqB8Jbsu0+tZjCvr7A76ROb6FjWS504KjpC9tGe2kxC
t/h2z2W+DrevSuMKAXHSbqWJYYyItKRBsctS3TfvsEU/7XSf6TYwGoY3YjmUVGh8
/ZFnaq15tkzzmZp/ZjiCod+0N4S11SkGxY+nLVJywvKJzfe0GZihyavK7UB+Z5Bd
fe4Zk/lJfGELcPneO3iG8PYi0y2T4aKMl5jBvG0ECbxj66+HecpPmNKlwnDb8EIV
bEKgH8k1y5hz6ydx7/ikjoFKtWuFdJcLkt2SlF5VVmMqiCAsLPUYHVWHvTJEQV+I
IefQPwXfXJ3LUNglFIa4X115LD3qkRa+80JBNMOW13sYYtWIorkD8tg+kL/lfjP3
Atvy3ScCLtjQ8lZsKVJGLg5nbDCAkYefi2bvzr+qvM0XWMhFyDpBv6SGTjURAlK8
Iq69qXMdlLDoinVz4/KaYrkRnQfAoRjYfufI0T1jzhlyp6p8hHtyfWBM0S/e7xtY
auvvZDoWF+05pHIG1uSZ+EzdAp7e3zptku2APW+LfpMa0kGvGIMjXbO5Yyom2IRX
e8l0b9RAX+azWzNmZsEiF3+1JzaQH1gRWcbeROptF6pZofBrpf/VIXnuYk/WYnNw
GiYoweo5+7LuxNz3aeU3ULwYqeotdUfKipz/dDsJH7J24NJnDYox6RB9ueFsPr+v
XetjB6UMAwTPyLcWiagHh7OQEectv53xcmwzQqy4aZRYgwrmOrrO9zeEmJL7xeUF
iZfFX4EQqfg+UX9PxPX79SWVZKdD3mIEVwFp4VaJ9LxaLyI2+R1U42XkC4PRUpLp
NDsX5t2Dmd8XOQeWlpENTaAOlsk9DPJSHCRRqOwnd/FfUTzzRFdCwyR85dayZX9r
BaaiIONdFI4vhvKbSh/tKVp/wPNHLnzVKTOcU+/z//nAbBzP5pEzhDKbpOY15XGw
lKPAwERAOdHFNOzdkS9ZuKAamKa8eOE+OWR09+CQFEIELFMim3sEA45I4Nprg+kO
FNe7CIrOzXF1fFKHQ9Larva36ZPpGgjUgiloKCpDCps/G3Ptpj91Ze+Iys3F7RAo
eVEKghMhBerFhYr2I/TBaop4yuLKZeen3ikSfyu6VoU8EJPE7W2a1rWk+XPVei9v
SqFKeEW6QQbXgShbTFkXFczRcVjbHYNxrzu93LnwAWV7otDbuwL1NDLJGlkpIKOm
bFPcr6tCHVr6SLXArnUPlK+HOYVN7py+m17MJCGRXyC+X+vwo8oFCufjRtQvvPBt
whnXVT99Seyu31l5Z4iRNEMxim1QnSFu/TsaSOWCX+B10MPwCB32PVO1h4xtCxiU
aAJ8tXAEn7m8SyV8GSSrjg3pPcUSt6odfsiWPnRQ3t0blVlkoxrKUhrBY4N9IoEW
lk+Rk+du38s6QfFadcXFqNI/EcjGHBB2ZXJsQusDZlZ+bxt1ydZMbr13GsSOMkR3
QQz22g82hR0DegPE/TECvkFEL09Yn4imd6q8dpjpD4R3FJGfWu5Fzq/gBbnYprw6
224IWgbx/uxHf2u9XQ+g8cTQcpzzZXQef6TgmaP7ioD2gn44LOgBY8F0aPDM53zP
AoXc0Ck/V2QsOEgjtKYRguHewcXG2E7ZNMN9xuXoYPu4dTrdOIsrSSjDYvj3/1XB
`pragma protect end_protected

`endif // `ifndef _VF_MBA_XACT_SV_


