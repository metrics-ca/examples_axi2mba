//----------------------------------------------------------------------
/**
 * @file vsl_perf.sv
 * @brief Defines VSL performance data class.
 *
 * This file contains the following VSL performance data related classes.
 * - VSL performance data class
 */
/*
 * Copyright (C) 2007-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_PERF_SV_
`define _VSL_PERF_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
oqQ8VEYx1w9OZAosvEgFu4kMbPmBIDwAGPo5jgmVBy9vqMB7l2ECB3liQbdOF8hc
kKExPcn7K8pw9j4yd5FZAD4A1DpmNIJEmGVUefdafdG9mDoS1MqyWSAzv2OH3gQM
RZhAlbNraC4o3IMTsbG8VO+L4ZYnpQdtVi+amki/90YLKi+u5l464EXo6KMm+O5j
k0XecOxI4JMnQnkMe+EUzmHCqDbpbyO6KWy9Li6WnOykI/Nq4AoX1eaN2UH8U9ff
7OlQYlErrLaTPQ5YiWvRkkH5K+wdW/w68QGExmL5HU1yyJUPR/0UVvHbUPACc1oC
m+jFR2PsffjHzC/PlPfXwA==
`pragma protect data_block
5uJQfHWqKnPTaZ0DXFT5kvC97rN0Eas1Ohv7nh73zI3jYtifQ9GlzRQDuHxnD/t/
/gwLbeGT33JLGj8OEzl+IbLfejgYpoBOzatn6fCmdXRdVvF0x3vCYp0rzdxlu1YE
OioT1nbYe0mh/wjDL7132oFPwqIPzXLLmsmekHo0PMARe9LDVNG5YCoFPedqVCjt
TC29rtCMCusIF5gQ7CF4rxAyDAVHjGaKhB3nTC6K1p3b6OnwMNOnlzB/VKfDmlMB
g2TvqSIyI4b75avMNfmEWOI/eqz9WpEmraXEroNJL+yPQKceUeKV1ldBkagdUBcm
8mPzD+4P5LsKOfQHAM7U4eMSHfY4Ay6LRAHkYkqocFUSpzIzaUQJ8YXplKnjuqjB
XpkHT6eWivaoofXffc875cb24zyOEHMtV46XLqVIo5czT7iPZHKGXs06shmRRXmW
KA/k7ep9zuUOGHddXHQPc4ytJznfWJd0d7HZ6hPXb+/FgUuKrvFz+ZDSaIfBOK0N
hcBfiY/Mj8mmvDDP8ltiiVIRNooCmvRNNs/zFB9B5dcQNMMqYPbKHJjpWk9DSHG9
sMke/nURFgy59+KooCT9bDLciCmadjBbwm94/PemvpRzbghfHo0ea40b8g+FNEhe
eE8nG6hhFBK9lXOVjaqPZ3VAUs/INJzJGRZliM5GeT4V/N19waZmSu3Bpad1O8q+
52yNJCILjWYTTthe82ewO2ybeYMIsa84dF5nIIZejFkTJc70Gk2EFHiOLhkkSb7O
iyQ7Y1pLlUXzqhd9yboH2eJiQIiDb0RSmlq9g+nIR1JFajFJGLjhxe4qXm53hrya
3VU/d5zrlCZLg8TKpMAeZ/kftNE15KhvcB42Ppt8dN+nC2XXfAfJLhWuq9Xpr7il
8vimsb+/XNnuN2vPlk88C3nIYnplmNzLiQIo9LrM5Hmr2QANnsRxAdrY9yKO5S4V
gY2bPqk1GcA0+OC03yt80wczR/gkDsDN4t/8cvSge7x5cmdLopzmFzCoq2LnY6R+
a3Rfdc/MBmBKgQkFHdJFHlM2+NfMLIPlSbMQr+0cDyc+YsJySP/qdPw1ziHdDfaU
/nNNofjEb8thRGw0tjrnJ81ol4+cOA6OKpVWm6l8JAP5VZJy6hxWD7ez0idKyMDb
2LVqO8zewsq7YALivzd6G4i6lkbVYqHtDwZnnCt4bvmXdD0PkMrUNtX1Et+cxSrs
IvOJYdSr6w1/+4ByewVnmvDe201E7T8grMsiuc44cnHVuPQz9bzc5Mk7FaaAraT9
opev4P6KhM5oJkmqxAvb4TIekq26dqaPekxzs8beQLK3Ao4HP9IdwLJ86Iemgymk
0Qld2d9i/08EYiDnOvvLwriqolQYpleVWtOzPXN+IZMKuf56TUaQ6vvMT+tbrAa6
TYmmFZu3AjFZUKT169Ty/euShC2sbu1CcpZtMNyS54+83wLUrNmFPN8YVBkCBXDL
oRPoPYHlM5cgnBuiZFGf2wMFmH4X4LPCrAQKXJW1RmuM4NHoSbj5XjHbFg9j8qI5
+2+JUUO4oOLzXWJhT/pnX5aVV4MtKN/3UGphreOI4rrfh7gV0PgEqidcUFJUwjTW
qFY30cPtrh1eBGHwrOIyZBARAoVJWXCiQgoBRnlwEZiYio/Zl/zOT6onY4+cgNrG
WVlg++mIilPeMU41IiCAxlRPfN8hr8FFjfD291YSUlPUjfS0ludDMGmzzwI8PzwE
qxC5Y9I246vQXJXNA54BfMvuGe/TNouQJZ+i6hsjHoBe6tNvpz15mgy33y4ikStQ
imOmCskcFVYnBSfehKUYNuv94Hs18xznUxw55OLK5nnXULJOG5sBY4kq/HDz8ZWo
Udt/7CvEuHZ4X+4blXb+k8cJQ8ZKQUXq3iytZQyCYgbZB9oYjiZBrLkz1WBiZJCS
6AEn+EQhwA1A1mouC4zHtsgpsaHXDovMT90AcgoHes4PqRkh72usvbvN9cqfHuDL
6hJuFvkmOyfxcx19ogdxK0voIJtt6d9gk8D9l6brquflwbRpBkSzJiN7eDB9TgaY
LkmBT7spOVjQWUFghHaa2NrrvW5iIJqeEf75X9W4gxuS5GbgVqfrN83kMMWUzBSi
HSHy07FsGojdNQ7s1N8MvpaL5yUsLO4yytE3M0lOp7Rd/mPQVqwnfXLVEZF+b1/v
5xBT0zqMd4vBf63SaVbEKYmFOnf7m6rL8cjnyUEGcuKTwHdG5aZE4KxxsON+X4Ky
LmzPO9OhxkMe7i3Sek9mkjamJOGaGVKnH2I5VtbG5bk0CZy5sELHObnCb+yMPyfd
Ao/271yyXAyRu66WJEBxlJPM03e+ZeDrSKLhegkbp2+s2/Mokp5CGvyPxSbU3Klf
ucPtTxXIG8NmJoeijU0FZwAiwQYKfphnFVSZIzBjLgx3tiSwBVJgBEkS3DmUDBZF
d+jI2zF0hq5jh+vytAJGxHxYdUkgcj7yusw8BdKl/Pa6Uf2n0eieQRpy7Y/U0TL7
GDiH7w26RPNa1ilLa0gnTpyPH2kGnCWT+j81Gt6fDfVPr1hVwVznCVOaHNC5HMUz
9zPeZLNbXwCnXS/+WFGGpmCiXFX+HusQVVcIaVaO1bYRlWmfNgW2L7RTZtiTWtW4
fuyq5PXRASs7Mba41PyoLtOlxIV0een6rtJ00ck037Mq9gODJdHMkIuh3tGIIpU9
6Yj7Ksbn8x+wlzKzFenyQ/B9TXHrwgH7YBy1RVxOBbFp2MLFocvs3/PH7lH7g94z
IOucJsmVBD3/hqB/SUfe6dWa+YMZEyV8LRjaplhGt6yYA/VuNFae8cPtjsD34e6D
m2nnMajla1ZYBXOfNQe2hkxyU1ozb9eyUyvNRJBeGQxr+u9y7RcLK+KBUkFfQ2lc
so371NSfpMWQPpyTeeR205/CfNxVoFOMWgfylvqQWKdBpDuueSbcfpBnRVFbdhNZ
GBcYbjNK2j7Z5WRrMrJdOKQu9iia6V9kB3ETQnqHr/Qn1h+9cr6N5Cg5S8WvDPWY
8LAnTODFk1GvRanFt/JH3nVw/KqMcEJ1tT6iuAQh/kd/++bKx8TgUZWQ8URFsi8d
tgWsJ/UW0PYF+5XggjZCLaJPcO3X2eVpTnKWFF2ukki3iq3Hmon7vbFlpahussmc
ULbt8xrqidEY8Ts9EelfpUUtUJ53oZk1m/jBscmk81ySLAfkhq6OQEG7A/CEPhnD
7GPpbSA9MypNRTQzL7nb/VWmA5vwTvYbDddbjZBK1QSc1NUy+raHDr08RNvV6/tn
qcDLnkH5RcBt1Kxe1ZrCeaMji4Sc2OWKTRNCxKeMM1uMy47vj1PcLrxeUdzLYi3j
YrPaA4A9ayl6mmQgLWKPVFq1AP+cxltdlmqKIhB/jPKjIWREuhMtZjbemhGbyU/a
15+IzETfLhFZqHsMjBNNCwlOMMiH2IsH0S6HNMuC8HrqJrom4IWz+2ejHHC05SS0
lOYrVjQ0T01kD1W1M32mgXMl6KOuyo9iQsIqlsk2gj9lEYsXbEWLxkLJYNt7Q4Vs
+Bk7rwe1RjgEhL2FGc8T2O+/vB9z9VE+2yBmlj2QBwoTTKtCD3EXcwguU5R6fmnj
GRyAo4gkECsPt3rglWm1kbL8Oo4nxpgOnoP3qXEC/2Lj3XTxHSOTIHuOUGyRywM9
1gObfWQkd+nRRL799DmxR1HNx4U0Y7DTLkVIPjMcOnaBPDvJHChBMfMyFaCfrAgD
SrJIDlwFKFt4O/v5d5pkwj/hxqBG6oU7gqGRgUoV7L/wM4b2E702iHpDwsRgj5QK
suLDs9eOFrWvn2jK1IafXT94YvRCfAlUMSQhk4GhW1eC+BU4xsJP9epvvFhxZvY8
vdaOmVKVSZ+65zJ0wqoADv9Q9Y2fRpXQwvuxH62VTL82yy8ZvhoqSaf12P16Lflo
zVKFbXK2EKRz4RfNquMBqP768+rOftq7oWVY5KF/hXzPmnGX7Ionp8j/txoc+aAi
GaCpjFufIYBrvMAGLKphXja4YeJzilySELVSUdUaZW/TlGCnPYg6VtfuixwJar8p
1W/VxZJR8iQofpkmHT5NPjK0pMN5sgoNGmLKpG0mPpvTDqa5KMPUS3YQ+Ms15n+9
9/X/UYVdUr/JcqF7XHluK/H50KSLEHI28yWs106uKmLthn4+YGQarcGPEaJDW7kb
gL4o3JrzxBL+SXIawPAXojOF6bQ7Bb/vYh3DDbTD3qDnBbc0RmBK9XE9dy0J76oE
HvJcGg71CfkbleDp2aKImieR4EJWhZddk9YKF96sHeTEDPC7slAZfvF/cbgssDN/
q8kWDIAb5u9WEApLRSRBW0HFkl21ouK0TvSu8myInC+EtrtRT5scIysJIIbyb2rP
5Y86o81TnsGv0MNWTrbcKcnwny93Dj7UiPsGcR8gPDVvKPMeU0kz1CDZ+z/cVdPV
2N8n6KZ+1aBctRLR/cn1y/w50or42eRGIuoOIwBMpYd3sCGoxFSpRAsyMHGkTuD2
D/323iIBLxcwh1EpJi051M0e/BrGKWjpDKxT8OtcEouFPHYMjFlwhWVHcxaol1p1
8GMEhQ7pQyU9Jb7BMNwB9EuScCbhL09tZ0QebtmsslI8FlDwZr0ThLS/FQ4BHJVU
spKc51EWkyc96PYB12ijMop6ysOCDrbv9nxPb0IHyn1dyNhZaLAWVRIsRLFKIKiF
5wOL0yt9ZzLRV52OZd6xfPAqaqNON4R7DED+GLx/RX0XFeg1RyFMyLgJAmXMcuc6
4Xyvjft/7Nj5dfPbcp121FoIfYytqomP/P+gmOWG+xCqQdow7Heu3axnS0N4hQYQ
aIMGR/dMVN7PymUbfx1DyKw37RNMJLpWyD8gc8Gchuwt8UIHDNrWoELWGz/UwWSt
YqZcBB4kkL6DO4J9i+NRBz7u54r8/QTRrEOuT5QLnfhu2+YY3aYbrMliY6rVD2gt
Gsha3sv1YDtWYOpBfu+nQ/MhjzhyGK5ogRP70g7A6cn2SHyOVshKrTdWmDWJ7JZ9
11F3SUlXpSzmPCehpyTda/qBFyGtP34y6Y6yqYUdnDfjuvCbEDyMLlx54TiJ8VrN
yDf085B27GXCUnqW3tvl5DkZgIWvWkqfzq9trrItdG43In422cL5J9mhWlxuyvSN
aHMK8EML4X5EKpmS/yfIR+d7LnMQcUbub/6b+O04cx8xumsiTNoxW7oYQaUR/2aY
TjNgaUh16EuKZDDY5VDBh8+jwyHCRpze0d7ZY8opoY4gZKR3r/58RbBAWPBA+lH4
XT+vQ1Q02e2ybufg04vVKR2sywgDGNMjS6ww8k4VN3Wws+iQ5I8YBOhggNtIZGa7
5mSwCAyZDrLwjT7UcoXYUho10FKAo2uPrqAlwP414vijT3HQBdD0m8dF/4X9i1hd
hLoWUcxEQtVtwnTe8ZTq1RddCH0jsMqLU+/CtnFsO4+NozpOGkBKfGvdN1g3lJh9
ld0/H8TDiYASL8Q/qoYXmETuLIKxNaF4BQq9Hd2wweuOPVS498WtQccTUHADDFzZ
50yY93Y16ToP8aV12F6NaSpLn+GirR0IoaCm5AYMwViSZABO0tzL5FOTx3tvB0rF
gyMDhLOSWV4jEZBWYJkt8QgNudn6XSHMTbbBh/cMPfBGQj2z3iAFKB1in8YIq95T
BgJkM70CGFEbbeG/7ZmengsvfeRbSDyzhRmEv2VQMoKodPMOYaVMvUvvSGwwTK+O
jzVPmOITW+f804yE6jhymAaS5htdmJ6AxzO8Ub8w7ziXwdi81RIFwg0jeT3cfDni
wDyoaaNUk2XU7qG08XBno/VVJZNz+YqPJ+pwLKJSQjRXmig+WvRMSoNl6Pe4L88C
Nl8cxAU2Z2jqHvrWCKe5TDLKP5R1BQmtwdJnzwE2uneEp1pKI6eaLyuy5XGwi1J/
/Yblcvv2YEBZ6bvQPxokHKGR5ArVzOofpD/9mIlcehxwrCN/l+BWkfRmS+Jf5Yfa
cqoDgoOCNLlOLAjRRI0Zds6MmDv562aumiB9W/QnHRS3dYnyEQdHZ53oQri/M4nW
85Z6HWUet7WHUgIVROTAG/mxOCzg7/gOatcGj+VUdjzkvAQLZRexc1tCqY0vFra/
dVm1n5dflZfE+w6wjQQLWs4bgISleRT6tVcCv/+Pt/L3lUFVBAsr7sEwUDov9Atm
f6XDq0XitLy606iGVUR0mX7y+nptoMIBUuOCpl4CAT/IXjQSvQDEEgj5QwnXs8hu
PgGlmBdKNfhw2C22WQZ4o7uuywurz5yHRy7m2pIxNgYYrWqolOgUZumjD1wkHr8e
0Z+nvMSrsG9pEY3eQ3LmL+01l83AeCKj3RA/hOPtcV8VGjdhLBQ2TgyUqskl7bDI
7OXD1xcAdnIDPaxRSNKOZ3LTUSFfNtXlazPUKvZ0nEdfTxLndXM9k3/ZU03koJpm
g/z4nf9MgxIde8Ndnm4qDzFIcpPq100Jawg7DOXKR4e30IrBwqkIS6dHSlS5PoBM
04hEAglHnGjLq54VJgY10jV+CDFVRrTk+5cXce1MhMoG6aG5nir2zgVu6Y7K/T3c
CRNpHIhPdWpzDauweWRk0uWzxxWPXuOpiK1LrTNdX4VESJll5OlQJ2Fi8t1XOcVP
xsbz8tF1Z++++SmwBtxGYf1P4RF0+TFdCe8ecJ+nA+QOe8xjuoFQQeavq+i9SlSf
JMKKsgXO3+6/+FRWmw9FpFXZ3onmHHDmHR2dMm38Q5DT0LIyNlg0ECLwmJFldnZY
XyymvKNcZKJbbjQ0n96/GH0EHdiZdmxfzBc+aSC3K+Wsq8DXBEvhpisEnCXRaXXx
45KTx8X1vp9lqRCn/qweqojIUruomKrnhgL52veV9SJ3NIBU3EvIAkPhSg4DE3L4
wJ97zs7G+wlDWaFsdjI6FX/kM+xnSrVh8b+S/9a7EhBiaCwC0ub9HhzxMMU3R+9a
fFhW4APp0wwI+TinQ0cDckmW6LjbVG2CNLVK7QeAjzFSKd5y9lfkHR+ZKFJOlmet
mCztR5Cy3OvbZbL9/+fFW0ZzLqHlvYrmeFIiyWrXevcT4KamNS1OyuXRlGRNlwWq
KA8R20FfuhyTLrt0YBCmFn+HrAbGKiRmM9wqgfSjcO2A12naDeE8bmW1lygYO8KU
TgrM7bcFTd4NG0vGHBwuO6ViXzRenx7On4Sr/ZILRsiEy8tRXw54OUDEX0bSBjQ+
0hFpLUo6uYML7AUoQanaP+YphM0FgCMYgXiRA6oQQKiDeSaaDqunOMJz3cTtu8Mz
mQjOFx1eCBsbN0vuKwJHOxKIpf9Uu6C0RUZfDOvh36TDL09VVQKZNe1EjcvX9CWr
zWeJC69Lf/TP9HFSWDDBORfiTAv0+AmS3ugA4VcDsVUHJjZRu6t/lc+o1/UqqcJh
85LhDUq5CmnxYJqLlVvKw6pnPeejqerES7UmOdoeXn7fiXrhXvDjLs7SgNa1Kbgg
rVnejMdxzl2/p2M4Q3B8YBJs1okjXKPY/PxeAY7lM+Vr6888eoBwYlKXD7i9RF3t
IN+3rMDLC/O5rktAe9C+B7uqQ/HLrF4nprmI9d1DzAKBvDzmmhuwvtvgA4KQy+wK
tBTZ1jhax+HbO0BQ1o5znsgcwyHgxoTWTFOrK+CO/mW9Q3rMRw5Epq4Z2YMpygq0
WWsgRtERxMk11/tfSBs77X5UaNSoTAo2azrH+h/mDTXTZY96qvecROPEuB2Z1xqY
4+D7EZ4X2G26XFr2Ri4EdU3AUiJ1zYvjvOtT98ATSti3adNwRHho2fJrSbPJx6JN
+O2WXyirOsmsaWlT04VCioVKYjsucX/Yl45NcJaaSM+rWOM4Y4ZdJUh/a8w22e7z
Ys6QhZqVzjhTb8ac+NE+0Ni1AN70NwjmX/GueZXxt0nY+fIQeQ6FdjcVqLiEHaBO
eNx3aD4AbNS0I/cy5wfgSPw/WGQP3VhoxWaTrAyedEJbxUyfCh1P3AqEYEXjuJHw
kbsnA/7oeXcbIFbJsDkdGuZUNI/cXhliOTxsk7cLsDwTvJmcr/s3WRYzgoqu3Q9h
4Io/utN7rcYUe1A5xp2QwmiatMGEjkBnDuxqK88guO5s4wgilyTfYFCeVn3CFqvq
/Rr1gmYmK1TFMqev5FDUN7wT8qky3jV45R9pGAskNoTAE7PtkRPSk5bk3tnqn3Vf
9G4r7EHIfjuNk4xtMUGaL6skcDxhqGSf9TvCCZeuFElAGErDbe8bNBJlcHSZdglD
fqrRBphj3p1DGdKC8Px6pC9mJciE4zbEqCEM5NR8jiCWBdTN8Ii904rW2pnrj2qw
eOLJtIK8wInOFX0rIxdurtII1RY84JlwvL6cN2UM4fNQf/3rVSQZej+oGRklYjl4
BQJlKxpcqpCO6wQQ6BXwXXHDy9+g/28Wj9i8OTxys9lTFWAtEqSwGywFLShZvHbd
eOJUwzFkRZVHSVG87idbI5HLSvUc+BnmJ+sds+ksKLxj0ZFl3rF5aC4LuMTrmxyc
X/2Rdk8vzgr0kK58QDvGd/swrFKO5ArRsIf+jRBDHgOaBDBiDQIUBjY/cHSnu+qS
yEtWQ3q+/53IlhrrNK7GAkCuDQySiyBr+0Rmn2IpL2y8AbZiP81MwJrBZk67VOhq
o0e1hrKdKz6oGm2SYfPF6JUiwq+UA7S9mWB3sRxj0/MQfSC/+yC/IWMpeqLIJjLV
1Gqf5aRe2snJrvSR+sjMlWHk7vdsnEFOzcsX1OpyldkXMspY/A09KFCl8d/7zetx
EFLATWCZhfmja89+bOFZNP8Cia1bDQ2zf3Mov4dWe4f/G75bFNA+a2LwrCtwm1ia
yLCaM9LyrcL+sJHFPy+gmc6TTwTzq4pru4c9JvCgtElwL5v+utgrpgBNYl/b0Jhx
S8W2PRk8RWYBSgZksPd1R7tuVBlqfci1M6kxN0ZCbK7mtu/ESLeLdEcT4g8Jc2yv
FZ1mvvsskghN+INj7Vfm7pnqsGt+ULT3W+LZTXiM1TZ69IfKoVYulVSryttWjcVn
K9AN+mWV1OoGCQ/p1EItES9XIFfOKM2NNtGAxfQ2c4sPLhLxL7KB1EF85/5ToVUF
U0X/+Zbl38TG/s9C5B0FlIMGMCTituO9H9lAb7Qm+QV0NV/6iGvqUI9DBzhAw1qd
Kds47PL0miXAKLtcPx3iGZxqJS7EZbzWTITgoE4m0wY/E+qGYT1YXDRIHXUoLJeP
aKnVAN5p1PzNrlzDt/VODCSfjt7ZVndu5Sa6BR1cggU/4rqJWarP1h3j+jByFsAQ
92ZsW9gi7ZSj0UvmeAmwYsDkXgsowGgHy9WbY7pKnpmdY5BgAH8ykepdUsIWNIGB
CMQJaNXQiD7P1vIcGd7S2yrmpI1VczAK4tn9NkZY7cu43TEEV2npMVdt4Xw7pOh1
5Et23e07700nvwPAPGsu77PiHlvesXI1+IDhcTdOt3zsN1IB0/jW2cGpOkhes+i2
LsEfwMnIL+ZYB4aHRtibzX7XEPbWsQ0Y9dSCTpf9072/air1KtGeU/dxw9EC8d03
9En54UdY4qiWNg3ABKmcNvx56c+rZ4ac7sH1u8V7zSX8GwJGmTOesUZBrT1Pan0z
QWkEwrt0ybYKoLpscPs4lfFDw6+lhzFq+AmBLQDwUENYd1AWDS4yXmYmPAhiEKPA
ZOpaEfmt9rhreKApCcoBXDkg562Nzf9BfVyOnPH3QK+BKwSMMrTenKaWKXkrOLoR
LPMRNTmoYH7ToapV+PgvWS6OP/RYjlHa9ZgSKAhi8b2mJY2gpiXIbRtuxyrgBdXa
ber8p1I+INtCY3jxwiPBU8TVUIfRNWIWeAxDs85mdTJqpAwvWkxUZ74wi/WuN4hH
LncsZBxDkvbmmRvY9qkr2i5aM2j6agsmrTrV38Ii1QYltSm0ZXtzBsyUkk85ttZp
/LbBDJOi1YhEKunaMBvd96LeJ0zgaIfGR+cSi9nSDVkTb2loOJ9ptvGrxeYJ2mER
gJG83549Djq4GvhVuOZ6aNzjHihA6iPgax0H3ZaoA8wjHrM7sZ/b912MuOBRuWuW
VRXhPwsqe+yXirw1CSCrW+loI7mB9k/cQ9uEy2+zEUZyWl9x0Bj5f6lffAmFo9IK
lznT92xzBpeimsl6lV8zrym2rzffva19LkJTXpjis40wJrc3TqV3XAhz19TmCtae
dlFC2zqMC8yldh4kNASy6akEv4T64TCGa0l63lrCSECh3qn/U/WFcf1cTxYANAg1
8l4xsuNEc0m0CEzFqpFXvR2ny0XhzelKxIg2LK9xtxw8IvLOpStYAIP5PI2TWdga
am8Wx0vR6fT/rO4j5Gs5T8DoHaiBLqB/vB4c0Y1EeFJCIWZDsOQIcgiCpR2RQJjE
mpAgO1eVamQ2uAIVj5CvBE2Lqv/QPRGdXyomti+I75OAuj151sp2x2VExuv15Bfc
PTY0bRCwb7LvHDmNX0EOpZjjIXA0uRNXQGpD6HDt8VCXv5Aau9tSsKJ07aQT0GL8
K9h5mMIfHtK/59DCD+xCSEVzkTwPysXBn/XQSX6f5D6ThDhjZMemCjrXel/Fvrwf
d/R3FdXKH+83WIJWRw3zaVlUujGx7ghtSyZW+zZ04oGmJ33KxFo1dZny5jh0T9y+
o7UIgddhfoyHmuFdO6LF5LQ1TKZPf73G8VwITpppiM9B+GXQRmeTG1I3gY2xzIHe
Y0XZSUBxoBqMPNouqBG44NakorwMqQyrd1x1yRbvc3pMbmtcdkUcqu/lYQU6JSO1
l42Z64OTp3s0EEc8Ye9bT2yMi1C5z8LLoOiPKnY2RlYUq8/u2MmlNcCsWeipYOfw
3uwb6ZpYbakW75LoXWuFSVJDzOxjTwFvLyCuY+73HkENXLuNtCN2EqjjQUX8L6+F
SSdVgvBx/wQBlhhe3NxlH479pzoXwcy4zSwhlC7MP2SjsUkPAWdAC2Oj2pNhQe+s
WcuBdnK+cSR3BOG0F/dbW7Z7YmM1yHMpgE1iBCqiXEhMjdVo0ymLH7EgIrXS4+IJ
5P7JOSuorT3ilYrhVJp7pcP2+gz9VLfh4DBNnKPdfUIrRozHWiavGajjhClSK/yw
+VZAFZAo/teHxVllm7qF0WBfi7s32sncLoredoXhct+GK6uLxSPVADOaWi5XB5Py
ZMtL84gU+86eHqQ6ClB7fuwof17ldCxE4e8Dyr2+uUnLXYQC0t7y0E0289hEfQ1N
QEP68IKhqO9xXEexzNji9kpw7UmJW9MotYtPc1R2WQfO1yXoiumARVA2KovZjmni
KftEy4xhf+rctjsvNFsieZe3vlw7TmMmd6tcJN2XpJX7mqjEtBq6rO176kSMHAoY
Cz7PRo5mwoTT+/lArPqMz2nlJV0/L09+9ofs8QZoSBAI9PQrfV5VrLHz8crVuZ7J
blQK6mb1RrVgJ8JoWLIOcAXuqipLWicYWp5qXVMjozxXSRriAa0J3ogPMRADYv3x
WoZFKHMIQZSsdUAucoZM7S3AnHU9JLmVUywkF2l77bU018cqFvaTraYRFdL2EYlg
0iGMplKWjR2oMZIP7Rj838+t4CBw01cRMV+7136OPmFXuHkeKzuUxHhFe3u/Z7CF
TtT2eatZ9nljsAtzm9XmKix6FUXDSMxBKOj3hrClzifeIvG215clBmKYBLvPoeEa
Q88Ju6351yUuRFSPTBoymnKVvjBIv63G1PfiDR9PKd3JcJL8yx3ZBQ6iglatAopk
IRPUQv9+0M2fzqKwTakd+O24H6mhrHgagGI3nr5cmF4HUf2zyvWJ5KQQyb3wQ4cK
ZXIlOgTh/Er7wDek9L9/8NaIJ2a7KqGoF0iRFVt9M8XMwcxzxjm6cGxvgtYC4eBe
rSA+UxGAt4Wczj1fRcbEyMfKbXID5A+r4DWVD9+Egc6Af6JnoQh4IF17PvG9v8Ad
abiS7INpm3iIWdUTYh9VJ1blAMUJSvgvopIZ1KTsLjHrJpnu4ULl4Ux80EQHlu5T
hmCXSw5qf7Gq45YeS/Z+oEo/1t/cHdpt9NyfM23vvyoVI+qPJuGfZuSJ21d/Qyuw
o6IxsIiSliH0IFaokGqwXZdOjY+MWPPt6HEiH78mdvzatN0pmgFAalVbQg+L0qUM
Klbr/e1LQuu8W0H6DMrle0s+EXEQD7gIG+rhy9n+C4w+FxJXNcuSfeKhQTnH6ZDp
/YTc7VvgLiG0NEy0l+X++Kr/n0EeLghCrtVXpRKCMOt5eVQqO+MXMs+zhfM30lt2
GHhuxTwLwUiAoR/iK+eBtWK93eq5FhAl2p3iFOgwa93x4sA/Ho65StF4AEqF+0ee
EzHgh18hkrIt0BMYaucnntPEyApMku0l/yGMXyE1tPogIOO67J450b9Dd4nNVEh+
CYCdzqzFKBXIupmP81+TthVzk0kkMfl7gtEV//noIILj4eXQU7WCzL25Jcgvmk9m
RSqd9J8Wjx65ax8qifFIM3EkGfCx38TDETvsb2bZ4x33Ma67cMgEfLxU4RQEWwej
hEOQzYfv/AUm6GoP85C2POR3xlmU+vRpk0aERTx1hOtdafUye0whpPtr5Bsy/DPB
6rh+LLISnS9zmbG6XVsYuUsb/eyEGYU9oq3iM/h3A+ah1ITSgAMmOraRoJCZIqqm
ZqV/8OBNEb3uim+2j6faynID3w8uXyNXPLSbsZaUQIrPDifzSTDnlDvLwurSvHBc
9BdD281K41ERCq0U3wHuMeD0zPwGacUsKo+Jj21lIG8qn3ihfFzvjrbqCbE5VO3V
3z1817GOOHm0q2fQspzYozly2rirIb23gPg5cUv5QsF+ECj7h944lxxzHA9jOfMb
jOUciRHvwoHhPTVb1oznsFxVK8xtLZHVAzBuvMCpRfXstjJWX620DFudNjkOxREG
eqWmgYw/LFS5zrOOSKOs09QYj0YH2oYVKo+XTAtctLVnknBQBKcU1l1AK0vD0+N5
wSqa2XHC3jmDc+Vp7l7HPoupvQQYLGG+irsmeUUuUf8hKTqypo/eZmEjBH0n1glo
i+NF7Xwo5uUrc56vVOfgT1GOnIyj8rcb9JSZKYzQ7/kHvUnjTa+cJhZ/zYXB3W4a
LBnasxBSbrCNuFZhXm4Qafx6n5LK6Va+zLJczo0cNBWqVKpM5d9wUEepXgQVWUAy
5JXKtdKNftW16KAa2KZviGXWhJCrvTT9koTR+p8Z1LfiPM+7/CaVzoIDefiRm31v
gM6rpug49GE+TLIcj2qqFNh5nio7n4tpNY2lq26QWtUTsX6x+FtZ1eGw7KAHKLFZ
0NQGkKKM0tYMVXleVe++FHEd+aEnIMvUPkd61m+Y6vCFN2Jt2Q765FY7f2h8K26x
8pFxNlBh2QfsabPUc8dJ4BBss2wlG3TyzH6PCkwD5lyEoXLBMC6OkknP8veNp3ht
HH/8CSQ6Q7Lcxj8qTczcPgtVW+gPuq7+U+MrPgXD3jfqSpvS0vRj+NQ3zVRFpCgE
IumoAIL4SUL3jzpXgR9UDXFnhQSum2fWyPr372K+NqoOxyp7UaQs62U91rlkgKlF
vq/pFk7ur+u5JCstcB8UnRiMePXGJWWaSEUc4FQLUVEJYLhQIF5W08EZ/l5i4a2N
WOgPl2dAbdPoTOue+dV4HGCfeJIGoTCq1YRzt8Weo9isENfhC03vzufWewOHtyDl
aR/V44TbtoFOfsKCqd5rv3KZocvLnYUxQexgPZdKMW/32TNVBDT1ELblpu30luDp
60akLaOzkKTNS9q1YmRjzaxwAHDGh7Keh7LEkq6jy89kbXAkehenDzkM7ioSWJAX
C8HnAAggYxIakjtrFlUf5PKhAGcEdaMrj4Z/UpiTI4ASuhgzsAtJ1PSN9Xto/AUj
PBK1gyP0H3SpIILsLKOkwulqwiTSSvFg7lm6JH9BRb2WjWYfvKfPP/DIp9vBfdv0
LGxqx5cD5KsER94PnBgEync8YtD8E7OV2DsIfnDSJxM6g9l+BtiaMIvuBYUCdKWj
kXExla9H84rU6UEr/TTj8oOpxOcx6bMyxEyX10YK0CNU2tA7BtConYAwYrgaEZzx
vLss7nR2Gy05oPkvK85PqiqEeHtyCti7XV6UIIH6zRrT11INQIhLnNunYOuWAUQS
xpey/xFshqXwkg5J8QZsQlHhNJZphl7PUAkc1gKU0R/rkN1E6BQdHd3AOfMV3uJ5
hZZIuLsJg19joSrgrJe1GKtjF8fJN6sZAd6WfdeWscn79G268CYCdPLP5yze3CNG
YOHcj7BnzZ10kdLLOtBKwQ+WMHZYEUK9q9X/gIrKvHCr9enMkUNVa7ZZi6GH5BRx
sg/Nw1ZuvTJylYwx4IKyEs/GFiGt58lq8ak9WkK6CH1opi7hDvEDgP9XN8DLIyEm
GoLe4oUQZXpio8J8j9bTqH1zXg0+Fpa+h77fFdbG/ppCpfPOdJlj5r+JCDetqf5p
NY8UWp0hqi/kMNkbRL44bBfaw8hvHOkyHSuoVkX+y392+Q+cEfjTaSreEMhEUTBU
/oXJgeuv2U7E3FFReKB4mYb0LuIDhj+WMGga48+1U2n91x3lqz9KW4OvITvPt3+a
NJ8JK4uEE7oEMnVxjdTvjUqly9Dt1r+Ey+v618xZXMhc/UtLBfBgtglHngZNu+Uq
uI0cB1UBWC4PfVXIYa1cw1KtGqGXbjpMfCxmBHhGVnCiEFTtGGIunrIFzPvWtNSl
PRWwNfRia5uY1mG7qdMQPXBayWfwGUGSkgHAchfpMRs3qpKjQLpFR87ZyRC+6+/N
FzZ3Hbk+XmQIwPltHNIRAJgI8dZtQoflZTJGX0Q903aMszQ3BiQLj7ojC8YlQjWz
5tA1b+4oIDhTdua6pul/scXuE6Aw5eyBvqEnxm6kuOWq848Uo0OQ8matLMrzgIGB
+n/k5Ie/FdNtm4wPSCyBpeNMAVkXByYc1Ox4okg0kD8C55KKRXsshMcOhpGBsJxT
27afJ3twbYzo4GDELkUdXqovtYVIZBcSHQGaXmGodcXoR8axKYAGRf+Vs3KbeH/q
2PJGIJhqdbfL6r1zmE/bA/G6zxqo0r8EbSHEa808u/9gdXs8ag+OfGeyAd6cFTsp
k6GkoUohMrNA9XfolNoC+b9te/WllXWj04f/qS8Hcsk7JsN8kP9FTma8mQ6nKQoq
YTWj0jeH8N+/sCY1Glj6cj1HJK5/42xWxlIJsLalGm5wHoNDaEAcd+toW4hBAdDJ
rgxy0pUgvK46likLLtwYgBpxOTDC7QWeq5sufzBYGDVGyCc1nMH5L9eXRycWffdY
9JEFwRIq4YSYtOh6CcnEdr0loCriqQzc/ycJ3kvwOiaMIYWu4p4bivvuuV60r7pK
gi4RxbeFjn6hJDa1IYZmVoLZWJZGGdN9rYdjy3iVxGHmxFevOZThUcWRVMhXLNO2
CFFXgQEcbeO0gyrshcGBmxMuVGA08EE0CneyFSEWBE09VATaXSqy2B1EMRSi4l1b
0i470hijklNdt9CLbZh+h/ZvtpAyaIFUlgLjbKAWfS8H9L6T0UY587z7A2tseSd8
CvqqYKIxDgT6Qqi8ZTI87Zu4/U/AAB51JuNu/E4HYWMPV9t7M7ZZ36OfDLwexR31
7iqPhtv+Kchf+TNXHbRJnYTGnKv1uBjO5kYADX04f2LH3hQfk6Ltb+AcES55Xs0d
w5J7zBv8iAK/7p3fzbLq5B7QL10ILEKAZKBJuvUDyp8//ZFj/d88tNLWXb9ptR6P
Q3Ovb3RBqJEET6EzBiO9YdIMIUOmSCRYv3hlxBlsXYiG8v7V9qynQdRdNRr5Yoeb
vvJ+LYpRfKeFAOJGAKd9lAcIeDIe+tfbpMdZGCdzX4Mx32JyPcAxy4EzxI9PYZJZ
doPjsII5Qc/h5kVplaN7uGnJPM/gqjiB0fHd1Finbyjqt8DGrIDpTYl5ko6qdD4w
nfSbdUjUpcBHIswzfOmDqxqBbw0uForkd4s88mMX2fZOi/ROKivDlkFUMX6M7UDb
V2B9yMlKOit7FK6PBWsn/eUm+B6F31FYcsnORwE5tetgYbUtcXIsvxgRal+n/wRj
MR0ff2muWSp89j/FKn/Zu/3UHH93APOv0buaQVWqCJTizKrSXBai8WAh+xV476tP
I/CyzEexZhjCIEcf5TPWEVdk0K9I/rEGeMJMYl2WCLPruJRi+wB0clIYHroE+XPD
SHTdfXcnFPN2J9yeTRbyqzxN8DYd0QzuETPLuGayB8Cjk6TDYVH8/5TsQm0mMDmL
Jbkg4ENE2vNPjJb7KaVvedUHzUJbtD6FEcJejD5feEyQt7QcuhShGRdfU5sf8v8i
J4HpWwyqm79b7ut89MNuwCjf0GJXWb4RsvmdoRCEyVo3EdUqgoUciaWyXCdpUHrv
cv4qJ/iURcBdGb9WJTL0rs1hML7Y7gTzVQhmKni1YE7mMjcKDlDY832ksmP8ZfSi
3awxOyjiE9KPlvqr9q/tyMR3bEDeV5THJwCBUinRGSl1GoNxaYLYJhEKLFfxx0gx
vlX7ltgx1MKEEfSI5I3C6neYLXjHve+Zn6gkiHuSkGBip0mmWoYT74JsiKDWHK7V
Vd4vws2y2XdiE5CTO7NfSMgKljyrBt+umFLpugMaehKTuBR0OwBalR8LjFuHlHtu
A13EsGxtiVs3z7/bAh9W/R74bf9X9joDxzF/D7TFFUZ82QVK2vnoBreM5vl4AUf6
2vVt/c2eRB5FghqSrEp2XbWo+i8NKp1GZTLtBlzUeHAXt3zthflpXJA2Z8jsDKOO
TWXalsB9zoYP1ke/kKKwwuS5tUzBeBc+5hyO3Lv5ZqoA+/ewZ3acRPifonKNJWJR
CGesqBdwOknuqiohR0GPHBBl9FUycFnOpvv6VX4hwJycCFf4mIRN+vFlFPoVnwSi
VjcD9OEiF7hWbQLoKpO9qhxNSaiLmy+dDZYx01stYpdvgFqAICbltiKM24eS12H7
AUSpaKq8B+HR0+0pn193IzjzN8xKpkOHyp0I9Lg8NjOiEwjLKuBQKeG42JlnGrR2
bV1TYtu2TarDuojTcyxwp6vgUCKWDHDffPL9yKucR09ORI/jJjiiiSZi8WBTo2//
TuNvpCt/sSdb50m1MTQTF6HQZ8Q/4jO+0GcLu7iu7zfMVSDDBNM0TOLIPTSEl0Sw
uL6Gmdhn2tSjxN9PmRtDNv72emC9Parf+W08Y+1Lo8ONqcPZ6WvHgwh08TuG0pls
KdKXUksEFdLgiW0KCu1XahCz8y9dl40hz7SdkLYElUwor5KyLJZYJfMZI53qTN9I
qWMkq47vPHCjUxE2zqZ3Z/HK7oItWGTXUbiiA2q0b/fXp8zsWBEwb+1GoMuFwXbG
KvurRTFpSRgXVK2CA5NtgqHorvAFU2b/DrAbP5zGptGHQXU/7umRBb2N1l1j4Lng
iaV+ibjz1lfXT9FRh1G9x3E7ZLFu8C9dbnn1xNRFfXwbmhlzD5eOre10TYNhj7uP
HfaFkqGCiAtgoC/vh0+Ikvp3+QcSivRMS0fmmC8EPsDRGwO+fe7pmLaXxg45JMHX
b0mRIfXpU0T0/uCRGmq7qipfAZrNdALJ9/gqz5AQmOzrl3nfFsBXeEla/CByIPse
XifSyPR5BzlNeIWg4EtPWqpukjG2zx+zc8zzngzaDZFcGNKt6ZuXZCWzgATt8MlN
riG9eVsqb+8c9nsseosDSXHL1oaX71Qh2wAVFqYyjTsikrXXPQfbCO4biWNSRnDh
OorquP0ba1dzICsiD6OS4AhBfMhZlbcNDABFaYiVPGbwy22Q/cYXZPzE5Ft9Pb1z
amMFfG2iVhQF2Uy4QEhj8ny+8pMi86y+ubxQh3eBYYZNHnFJygiJ8zL4R1pBh98L
SLxCpZRK/Qy5onO6IHjKHtq1LzK9cH1QJi+YVyvm2Z9vC5SC5t025UquN+Ml+Bih
EVk+5PUBn+O55PYpVSntg+WkEw1EQKpL6OFKE9VwkzAN0TNhXr19N33ZafqxYeXG
BtdvD9w5S6bArwVo4WWsC08NG/bDUy76VpAxHJWgv4stYiqdJPEZPaC+1CMa3i4l
EHV9xHyMPMTN+VYmbZqONadD7lH+6AlDYA9n98JLH+j+2I5VxWa+VU7HuVwwmWU6
bVeH+Fj5x9O2bKLSAISakk+o1I8LOY357Pyo66ouyrW8H6fuy7YfNayAQS5jkfUy
TYJnBZdNMFoXdAC75rw85w==
`pragma protect end_protected

`endif // `ifndef _VSL_PERF_SV_


