//----------------------------------------------------------------------
/**
 * @file vsl_msb.sv
 * @brief Defines VSL Memory Scoreboard class.
 *
 * This file contains the following VSL memory scoreboard related classes.
 * - VSL memory scoreboard class
 */
/*
 * Copyright (C) 2012 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_MSB_SV_
`define _VSL_MSB_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
GW5p/FKwZ+fQk4kTPp043TeRRIFSUbn5DS60EkpyraiaAMVjQc06tjHR+EbKfKZu
Vc09LhTB7rSyg0OaB5dnGxdlx9rQ/YQ4k+P8xYhzXOyyOtZmq5m+HwEicewVXaiw
2y4V4h6UNocZRe6c5tmgulxebNIFAw5P/ERE2fuakfsJ75FeUfM6V00OhWirUN0j
W5L2/Wqq02zWAX7DsXbewlFAndDNjqolGzlDfCD1Yaq5n4eOaMnKmYvrnTniso8R
PP4oAeYgc8wzQhdpwFpe2rkPdBdngQSrE1Rr0vdBw975hyZYlU0Yozgx6XOSDrMA
Eq1KA99JIfTdHiDLV+YsaA==
`pragma protect data_block
oL1p1gK+UQrKmXYMVJfUWi9hmXBPay/oEHCMOc7Ww1mWy4TEc+oTBJi4lLQz4leA
d6qFiSRCTBZXKqfAeLWvB3UDLDex5ZcqGWxBeJB6YutUTJEueZ3StVFcwi/0ZFti
txZKBcCxvumVh0b/9Eyb836+Yp/LwO5fpBgm0EHDnzJfgqHPSSDCJEkJH96Uu/jC
+CsBqFKH/mZjVIKcJ5bzJyJxM+YTeCCuw7EzbkpLsfxvBoJeyptLgKNHu6c7exXa
rpjPiT3eaL3h+P4HYXcLjrSqF8tSMktTcezKpCEP9o2PE2Sj9FLbUQ2ftdN8qypq
9ha5rrN1eXWeNwWe/P7aKyGEVAvINGnuYdOJ7Ekdc2L+EvSDKbdKoMgMqdGhlf2p
Ic2AqTXfCnnH2nsmnWUmTva3HTA+ZcrL+NQEre0lSs5HHb8tAEVPaUYnHqOj9xnI
G0+zpu2v4tx+mdSGqIBKoHfZ0peOOM1JpEQarDJy1IM/2fqTSEunMwr8ffeH1HAZ
u812dnRSHJscnWrxv58IzBHTFfcsEcMJ3yFwN26CemgDdvc2UN3vHG5LGVzcliPh
2KFRbiZwB3EqnKj1kJVfUqiCK8n+5Q0yTHbbD3e34w9u/Mj5bbMpiNzH5rjYnS5g
2tSuLpXoneqJrfkmvA3hf33xdHfZTHA/4F1zmkl9B12AHIarZAYdez5b4KIhWkd/
2lZVS4uB1gKgjSI+dmjkeKNFd4PBmBkWI/vwmZQ7/Tuy9K3WmVLJEfAxOBM4l1Ke
BuYbkvvsNolj2CrvqjQt2iWud+M9XxI/WIP+YTw+5nta8C2760j3b+gtTUMrG63J
wpvSqD45tuF/4NFjgnXV73SoLkeP6UtYViG2rM/ITdb17nhArif5DGjoFJmJJq7G
qBQVjnidK7oqVFxfAIqJh2lfi/otJLgNhsO4BGNO1yMxsI92Ap27sRHIwbjul3ab
GEsFXpl626wgP/q4D09dW2bELgqjqXA5l56uW85H1DKpWF5iBu3f6dG4MFr0/Pmu
z22+iFqQ1uoQMhxdYdizZJ3C3nEuG7JDN6BMLSZ7vlA0bw+zTZmT3EQIKE1Zsyds
hY4rAJVrumcVmsoBgGKqBrEyjIUb1gSEX39ZtEXEQ8R4/QfyTJ4AVDvH+l7YHvvK
P3LRhlsTnb3Q0laqLeg2YIluTNyFSyfBUrgi65bcQy3sHhkxgSnzbuoo7fxgMcY9
js0CvpKorpG74JBYpk6fA+OzE14pEu2ir4znLTV8J7CHiYp2pcN66MaTUgi1GUuY
s9J5AMqHi7OwwtcTpFT0wEeHLV4CnpB7Rh1YE8hh7cgOt/LpL80b/U/ILnk3rOro
H5K0R5FdGXRaSz4AKaQFgD66aZssao+1Gvo4M4qDC39v2mxAIuH1ZSuiboIYO8Y3
ec8ognzxE951sGOzNPeq6PKWIKBpZv6KFY7ege3liHMzdoKHNtvEZvA8cpc86Pyi
NJgp/Pz26GfiQRUs1WdGGQDAX7b8qdBuHpX4cvoWrEq49tAA+48ROgKmypE47bYE
TVJzH8wM4zsa5d7tiT31tm/z3ZLR8W/PnsgI5MuZGgC/6rsLNBtSeftbcKysZhBD
8NeH2YP5s5pzF9aAUc2yCC1zt37/H4GrhPMwR7PGPvyEge+nSFx//uNV6L5mmTyb
0I1GToogcyATfrkBi2XCHXGMUy9/oUKuSFCLvC+ycWy7i2an4QyxJRVntqdiRIz2
DcwigxX+W9KUrRqd4zOxLJypH+D6yr17am9hyGMgPajW4k8px6x2gF1Bpoi6wUv5
WzmaSRKH6lbWWdyKRfoHUot4T28R2z/2zt+0URzXaU6ENidkaEmqxg1haZjS0hD9
l0kBI9fcwA18UqQLDrV/04A7IFU4nBWHBF8zMGHk8Iasub39Up2Wb8+OumpKSCvf
R+jMleaCaJ0jVyFluWR+65Waq9j7/tfAOtqaTMXP2LC/ZqJkhbgCJ++D79qY5HTO
ET3YzvJaKLNi2D43aOmAMRv9GjDK989q/IUv1gTIWa/IO+Hn89YzPUEV7S+go9d5
JVYVQXOyuhhzGWGF+FRb5V36w2zL/AD5fOjw4eKYrNlx1w8bFJZ7xdfUsbUS1dJN
hkTe5DUsBORioWWbm+ad84H37jbHPGf3WJiHZQkycISdBrzwJz3cQVpgqXqCWuCJ
cxcmwt0e0pQb1xORkmcQQkil/ze8F+8JNU/XZbOPnGK8pjec/v9920CPcc4ek9p0
Q8Six+GlSnbc1ExvKoIRf6BtUwabnXx+55k41/5EbN8YQj2uvGyzeoj6NfeD4NK3
anEEkgQjlH6NDtzMgty1ZJb8aqlQ8jik2tA0opldwWsoo3z7iHCm/y1e35vxnAtL
knyD9t6iFZUn52GU+tW8cZuk1jisbWudWw7Zj5rkIifuO5hgECjp0K5u3pLTbRbe
lt5saPzO9TNWBMUQs9sHFpJ9zh5GLvgu52j/lmb0GUh2KQU+rNWiOthIy5KXR/Qb
7zCAy4LDZBLEbvgawjb7uUi2zxO7vYL9yqU82GtxaiZwKMKqZNmb5seokAS6e34z
jt6uj7dSiszLMwH0B6QIOGqMs1GbF3TxnqofqrME1aNV3Gu+WuOoNSBowgGwJ17s
Ws29AqQeqFELGTotS8ZeiCVXSZwc7sDWO32btOBd5XT7+fAW3Ua9m33FEi4tHztj
VAJIfU0aegkXqw/bGoLYmB9y3+fAMp1DNNPrVi62GKz3d5wUUlcAcJ1x66E8kRHI
L9mnQdRxoKeR3+iGo3XYQcsWFN8E62hTu5oFDg2g3P6gTc1BLcET9ewMlC8kcsJS
U5TDyzDS399BcYH8is680DlJwm8ZVv6seImc1uIqHTdApMEbiFaLQbh9eT9QVcsg
Gi3tq0shiLeN88DUvecZ2WG7LSHuSxmO03tWa0ALgAdUuGvQ8UCbUDJfCzrkho6W
XD66ih0oLZ9dY1Nz3ksyer3C7a+55Wb3K/L8ayJD88UEs53K+ji+OtDeezTLLzV7
/H/V5mrS1J+Z8b4wWEq+TPNFdaWAX8qKq4AGf3tTrprmnzknRNpyC7kdFKDwvXAW
Xvv9aPD8cew6nqlc4DNNqsdmKi7TfpVk8E8iZ3nzl8Tse4r9V9iENPbpBuWup21R
g28wUza1Rb5OJ6o0bDf/cHYYjB1Qu0h3KuNgszqKv7EnDyrxbyWqJBP7eq59TykX
8Rl38+SdBCDLU5x4TBv02JzBUb9rdLLaHPG/fben5nlq93Y/eRp0YR+pBXPHYHUu
ynfpYmX8A8P5cNyZ1lTTo7nGnMHX9tU6U8cisg1b2Kg5NT8szET/JrLOJv9cbsKl
Bk8Ejt7RPd5RYno6Ui7NoO3Q3l3P/fKWq9go2D8qOXbiJD/3ZdQCTypp1eMdf909
R81wnTqQnVEdvOOGeafDFLvusdNZQdEALgm9F8xNkvS/jqBqH/kV+Vc/Qkcm56rR
S7P9ZhxBGscgdYTWWrG4wyThpYvVC4BcOVqnFAu6ga6OKohMyxfBfO1xK/aBHx+C
It4n7lPyjoA0nmIv9bImyhQa+jeuBgmX20OKfp5KpfsbfzM877V+awLwvLB6Esz/
fP9pYEyWql4xoTCYSN8jnvZkL6Ql5YolZwtc7ZqbXXBUWgHOm4oCrMLApskZFqMX
1rYICr/m06Os5n7yLLNrCPOO2i9qh92xixYvl12yYQ2pCCTlJCXGDTOP2ZKwFDIU
uQJhD1qEay3A+EFfOYVaUo8YCEbkWEqiMM8fDCwWyMBqJGwAKHm4J2KGV8qAQmeC
wsI8oOaaozJ2hHOJo0wIzwsmtlCmQa397P13bk8val6Kk9PUWTt8G+rkeAsvBdxO
s8ShuluFzQUl52uUSjh5PfM+pB1WQ1HTPKIk6l92XwewUUkz3J/5Sbl5V5FprFt4
TsFNwITKxYIt5Hpz07GtVOEiZzbMCk5JYjGmaNaIHyQNwk1gkdo64fXTuPs/YIrE
JkWk8vFLUYjTLsccKWaKpt00GcK0kP5czbuGFPwFuoOnWPg/PqcioPvBD7ffunnY
Q+YC8gEziQU2lLXpZ/caePirkZ/Sc4AWmlh4gKjMa0KlaBZ9sXGWFofZoVGNCxb5
fKvDzWlT1U+EIUB9fMqIagkQSNJ55BQWhOh0HfuDijJS+DkFbQBAvvh1WCfyiPD5
I6WQofMZLaXg2l/FZjOjYQauSXkBteDHqNMBw/awbgv0aczMImNFBZz55BQYFWLM
Y6w9HEMmJa37Qlv7CSgrRS7fWpxllt4oK6tHolHMlpKj2Q3VmPFQXiZ5+J3FHVf7
maD7QxYUthWF1ZDm8AAMcm7Hv5dvZw/mSV81Ses/oTfgC+pKjOsjbs0P+DJwuvrC
K6bqzmM7+KC2CcCzQuynCz4TW4PehXVCBqsbV/oIzSiiKLAMt+ctK20AnK+Q6d8k
P/px9LoimnT0uFhYhckm5VrXeDXpH0DwBNn9rLu6DL86O5mphcg7m3XO9SC8GFIM
d9x4+aYH3kqew4Gr1fvN9P8LFDwvU8JXngC1uDp3YFYhfHULvVu7Edrqhs++hIaJ
70nlk4gQ7VhoTHTMg7S1EIbEV+yS0mz5ms5FfeGOY2ikNw95XovP+EtGX5a5G3zm
BTpH1wp34dprqxvn14qstpuw6lJ1E2guVEbXmoFKDf3ZU8DnNzHpl378rvsC65AP
TmkrRRGeGnBa08IH7523sX8i7WKMMpZaxREE/GE0KKO61IyA9wmeZa+Zp6r1OqGm
frK1l8CW14rU97Ee5/Lye/+UnAR0iY5FOrzeEOOpJUrnAZYyooDcQhRlW3G9LIfU
jVfxpuOsNtkODeVduUvrPaPEuM1sOtREGHgwC1JmFz8uxfLBvh1Vz/J/HMJtW7PG
IzleVDR/jptI29tEc8gyJ0INWeo0pV6hfd/ODxrMyA21HG/KIb7KU1eE1W6p2LlN
RZNG7smvT5+f12ECGw5oPokGWeH1jeWqP2wo9+sOUo4r9wpzZCAFbKDSoq7UYs8G
juvniHqPuiKh2itQvSq0/amVyhN96WraCCcoxj61rHyTbVWtuAEB3dEv0P6wxzNn
jrkgutu4QrzKb6xEDa9ceSHrugzA6my9iOXOvF8Q/DWfnRijApNZiGQB80mUtbDQ
9LeMJ5tFn4uD8Hi6nRP9DkWnDoUn3xMcdrg1mioQf0KBPZToElwGlAcu43iyvqnF
izZ5s0jIIQgU8IFq3BIqg6mkGoaa9oxQaQM1WI3gZIGxtPwfrPF8fRg4bcnp2YSp
vilWHrQQUvAJCpAiSiCwLvxg/xlyTv0FxhwLcBIAFjn6AfXMuZ6cK9E4G4jHwlSg
Lsw1zL+rAte9kiPKGca2IJi7Y2heRpFOYhlbJ1GUKHmtvM3AMkju+OlhrslNbv5e
DMBnYDSyVxkdzg1xULQearMyQ0c/mxk0yXquGBZdI0xnme0RsA7mPxOaAipEztV7
9falhrx5QHZrLnXyI1ClB3RlntxQHgkYBO0lU4RfgB5RxU6Y8++HWpwz391RUgp6
m46SmyJo7qobu967XZ29DP4V4rxCKMnmgCg99WeT6NAPfJ2/wVFQaHvCSz6EM0gK
kawKxaN6tIeFHJPFLaHC8omQ6wE5o2npL443Pdm7CXM+Qr5G5edMPDHA7cPP0nMO
g5PWO/vXp6qR5XSET0nvB+tXwQANVND0DUdjJqO7dJoCX+dbRMHbs5FTZbwvNkdk
p/n0Yo4mhCfXPhaJk5XohPkxZdFtbOFtTfCp1Ci0c8r+cw0txR5AyeHY9O41YkbU
Y++CoNi4J0K6f75WpySL0n3UENSgja4g2y873lLF99Rlxw4seAnGcor6n3YxOtnS
cxybcndVX0CtmBkot2Qo6ampXtLpS/yHYvJRJ0c82Zpmcu2zK02mPt/YAZv8xHHz
5SVkaZfqdnJEnb3GTVGZ83tjwD50FiB590SEdV/LLMoj/1+a4t60t/ZJVYOqAYu6
Vh/B30icTECbrHjDHgckJdpCVufw8ymXzuZjERUZX5nW2gy/CmRAUeFamewT5J3a
JWR7ebYZBW9utP3Mt2/Nt2lmcT+3XdA17lbXsPD/FEHh59l6zHGWdukSXPuY1dvZ
MkFYfNb4NYRkpxQnMi30foXoyFPAuv+3kYVvh2S9F296UsgtVNCNz7C9Nhqhsi2y
KsUqmT34LuNYn0i3ng2GaZsyyZTHZciVHUzaZJM0MnwdUUkoDuA9Riw8ctImfmIF
Vq5KGpRxF4byMfLZnDt/58NQAwXbudE4BToKMu2VOD0orVheoG5eC5bxtpNRAZ5H
vbvigfgvrak5DkVENhIOHh2oqPofwgIGDDePvTnxVWqaZnhEG7RvXSRf9ahrmJFM
UmpwkPG3wQBRt2PdclIBF6ScyrgqhWAmUXrWBTX/9H9gxpaWZFPS9d5RYIQKK27W
BCn6nwV0Ec1hOhR0A5VTZXLBimP/jA4j26bWYlOogUkL/ATzQ1yBqWT8vf7axCWV
u2cJ8n72RUBl45Srj/8PHIZsHFttqwD4fOYyPHu+wGsoSF575ky5pAsumNEP5UNC
wis+pJF0DmChDchvJqWDCmgWf1uIyqk1kLRpcDx4IvHXrXxse4qrYBVtYkAQgP6W
d1cTkOXDrPoGbfZVFRmNs6dvXPkr9y9mMLqtPK47JPMNzdLWXATbaIonibwY1Nrt
X8QY0b8TsHmtf1JgS228rIdT+J+lkTQ8+TE35fP9zPyYBgSZ6DtzvFTuwTy9ElKT
oQtX1b2VhAA7517ItJmVkFKM1wUeOt9/f5Vzpo8S/00N/u/Iu9ZjpuPTptuelx0F
hKiFXrgbBgECagDsCuqGLRD7GWsIb14BSOZiyOEb5mcajNndYdAAuTVAolMr1xqt
EFKDyGXJxMV+T1mUmbjFI6LzaIYDhFzEm/ittPhw7MbZDk4QWcI/GitPdvu2mGW0
ArzQySHSgiEEqmrqNBeqgsosfXIFcAeZQnamPbJA9+6eLGu7lT2/peqaOQKPVNIy
Oukcc4F24Pt2VLWwgc7v+VbkqUQk9nsXpE1HzvSJlzwYl7TPb2zDZzvyhT6+PAup
7mnrKKdKa5odO3mr8ldSQncqsgjOSCmqz18UOwppAB4c9L1cwmDeHkrrPJVTattm
3FOW2hNaMDBatGbU3npQwQVl/W6v3kJ12+WY/9UwF541QEA0QQWhXsU+CtW4w2Us
AgB1U6OxgtqOvAIyc4ttXC6vy+E0P7C27WVniNbMGaPL2EUjGo3UajXICQXZVoCT
upqmf846OXbQqS3tbP3nH7qFuZIgLfmeuUrlsOnk15KacwDey0Fh0rV0KLD0gTri
PgPKlz6L/tITv4pmpfZBvfkUHjIdrJYMcUDJTyJYrVggbZJwG5QA38QFr5RSlGE8
j3BqCyAGkGCnen1Dn+Dy4cM7r/FEXdnhfeRFQUT8sqwYqO/ux1+jYH0D08lHqvnj
aegqtixL4WWQ7Zq1P4fErkmwZDv0w0MSRdJuoSJ49W+v4t0ARldluZi+Hhgg/ixB
jSicYuvsHxsiH/jIUzFeyKlFiUkjDCTuBP2pkBG5js1a8ovnch1nte4DJ8cO6arR
xSAY5FjU79CZo/oomkGVQ64C+ZT3AZNAY9JurOtheCprvbnGVblMkvAbhyl9GxcC
iiSIigP+X2C8ZAaGXczg2LHVjnKkTj7UcFW1rjLJnm66hUEk9OI+B/XOGG/b5dyw
ADAa32x7OHJ3FSSZB7uIwBBGDswlmgSG8Wwx1ZX7K4WBTeaYvgLcwCAQjK7Qq3K+
+bpN6AvqJrTE2iPq5HCKQt1vF2bFRrqqK1j1LVIVz9ClLg0RfSF1e7sFspGI65ML
TPKh4NVyfeyu0jj277vQcOjdRh00+EW5Xk8rumHuICnGhq1EjfQK/vAdiIgegp4i
ECiYd8hY7X0uTXf45rZuqPR/vJhE8+FOYZkOC9o815N/qZIUTWXgZE6id9OS9Qq2
LyTn7qAGovftsGnjQ8jyJGbh4UVKopYYGvvSEjh514VtJeACmIakk8qQtfnqoO+B
5dBMna1xAR6pGSQRyk4WUy9ZGveuh3synifATAs58NxVtGVrlLIaXXgCpFBUAJOQ
0cwv6DIvYuqeWnj0POm3PSzXvhP+lJwLZ+dm1d93gLkdQvG8Wqw4xQ2O7RqATQn8
sKXYiv19tJlFjUs++Dszy65e1ysEdFXRHVsiHhVy4uomFjToh/+KS6jvMugDSprZ
uny9gGGx5kFA//b9e1phoYVcA4wvAnmFIfBdqVyBVZjOmH6bQv18mEc+WG4M306b
1h+zZoBQYic4mh3E0rQsZidzgUc4TB4ODQSJnguStuw5ND4deI8vRK6bTGTgvRC+
ZiBojzPOdWUu3v71MVQL+TWybznKsJHrULvwiboyDnINSMpO5eGACZ76qCqI/mkx
0TZ6B7ZRb/rqpG2+Tz7mcE9zY6vW+U+jrhZi6r82YdTYWs1svq6YfS+Ax2swEHLV
mlTf6o8z2v14ebc0NNFjEIPdw2Kif++3+G9+oVghHooJeQ4rVjne76fDXYlKRlbg
XjCECABbFgdv1qszw9wDCfmc1vv38lETYrZg6TnFQXgg77vkhSwRr+b+JjRuU1q0
NmGx8Gg64ytY6IEwAy9hE1m6dXDQcuGqsaKStYYHQOHEPkfIAVYvzTXNyIP2Nhtm
Icacy54jmSduALz4e4n8oI/hyqCmHPMzXFvTRaGDQkZQHWWkQ0zZQBhoTYcr/tPS
qCdRPiJ+WJHAvrW6AFWxDBVdDXJP7BAmBVZRvqEKFXMdlNxyFn/7DZARfj7qVQV2
xEPBQZoTV5D0dSSTrKfuRdWW3bACsqraK2i06iItXa9MBMhuDvkM+38gNnH7pALc
2EhuiaW80rXDy6FNm+ncJgyRc/GdzuY1sJDhwcu2erBGhZWkEVuI+TCXMZH0YFSX
KXCddInByPkvucxRXwhIGI1xY9Rx3oBSa2xuM6OQny/1S9FiF0FipUnpX57AE9pm
02mh3p/1le3Cc2lR5ssDAdMNslpT1JGuI1WOb5mnHLad+W9OGkcP+jVNrwCgxVNF
+pR7KISVnKpYw0UootN7wnXP82GRp7HnAp3Pd6PsLC2r3W3tMD/l//B0XNe7KhKN
ONIc9qqTYGkSN+9rYS5PZOg+AvFS4YcbGlZW6i5Xlo6oCXN5fYn0VgPm/L0rIP4h
taQYpVpBzASsDfBWI0G4BvlwfZEAfVv60rcRZCxISV/9bKs0yI/ef/n+6HpiyWa9
bZqASpI42/IfKzjotBB7fBg6FaNRpTm3TNPBkbNvxu2+l5yzT+sSBrFFmYJzyN91
SDLuI+NEZVZjnp/eUTk/bLAoC+lUVOsOn88XPzZXnNkKchw6UIV32qQrJnvviS7Y
nhkfqF/C7VznoDo8bgR3drf2dy2fJUvQIxjLZ3sisay3H/f47Q98byZq+jgJm/ke
F4j8hEGCqh2xLXyJjk0//N70Rz/iYsQ+Lt7XYAg6zOB1wZvkyT0utnDFbqnSRbX2
mkt4Y5Vvj7J/c1JskIhr06xRnLEiwcdwpW6VflWRTOvd5MYooaOAb1K5jwPwVUYA
4Sdd6g4cMxtEiCdCuXoZgJfDQEA/dRw/qS21PNWplXa136KRvdL9m2dM0IOeXoPP
qsxSB7O+AtfVrgM7IwudBYqU+3qCn8FQM52IaSXxSl+mUY8lZ73gwCdROgieLANI
9bgPlhsrsTPS6WvBosgYeo0nWzlM7TGxoPRNFDHXeJUafjwnYFr0NBydAMJZ81SH
qqrtmjzk5QGJU7IZOwLvZWWtBYXs8UYUUpZLZZ+8Z7gTKrIPfXb8YD3sj9ZTtyd2
MT/ZSBRXKkhAtCRtAceoAP5LbWsYwXOyt/BXM0BFKzBZq7RpP8zi9EKRuTp5dfV3
tJY93Owdu2+Wu7LxETgwkA/cCOllGiCi+mMK7eW2OSNh2mEeCjFZrRnjppb1jdc6
APm8ZJn3u7sO6cS629nsHyLzlX8uYRRb4wkWdmn9v3XbpsCAxPQYJliPJKkeubrX
f5ao/f35x9OxeXwRVrlwZdrms0wBpeWNNKQckwr/WyDQPts5BZhb2LbSdDlZl+M/
D/mwoSEC7m0x2KglFg2od3qRd3UE/3Ws+yQFkQqn3ySa/QbwVH9j4c/ru4nF/VWX
gTNcA9FxtlEiz5+FF5xtDhgM9TwHuTVd3PCWbs3O6Va6+H6AGhYLWdveBXJDuK80
fxdhGHCo7owPUZBUJGLyQtW/LAH0ACHouXZRhICnpVMrCn5UXbCKn5Goj1BS3i/g
60+ps2NbiW83cEKHl61NAM9E8MJZIU8VdWZfQgXBVJ/zotsTsdr2hIW/kjtqqft7
PYYZjKmq+y5fSn3gXmEfGeD7vPUyIOBGqiicqqzhOU9ARou5ofSLMjeNoA36Udq4
7brI1Oymo4M/aIdIEVgP1C6+Sf9dBQcuUDhfo8xnWU7wR6sFK6JghbieI6f6NPOR
N8BlI6v9ADX4uThjHGk9Y/SiHfRllit0F6qJJJdsN/4rvCYma1J3aLabaG9leUEK
Qo2/gp4Z5PytUYorOW5QLuOdMMBaVxejB21BF+3xrz5Wu2vsAUHDsBvtZmvKR8Jn
EOoaSozTVkJQjHq1KvQo+Z+LjzFUc40zHPf65PbTWu/+SB20iqHUsmHt1UC9+as/
j3rl6Z4U7OObb7qWmPQFodlLZKnfJlQBwGqzWbRd6xFFC+HzFxMF38Fd+PZbbglB
TmA0xpk6MVNRzFQlQNQOnSp58Ou0tYIxUVkKTR03gfdIfhCrIoMqekpYoH2G73GG
aaBfdDQIEIWyQERr4DpbxHN3OyQO1iRta5mLvLkRvC2+3R+j3OltJ8xtnEVN1w1g
f983NHSfLr2U0rpk9w23dnzGOrZ5QIsAZPuNKtkenMSaB82tRsuCvNIT5iUnPAFs
GNgxUtd/zTMKLdvdTybFn1/WncxesH5EOWWxI6hrzcHUD96HJif1iuk9KSDROxkH
FKdfZKGYa6Dop/+XZ2zmZZgJE4E8C8rl1qjA3eDq6oVCs7Vq9VKXJPJKDIQiudws
XaeYhPmXoPAbA1Hs+EimlCl55LC7T5JXg7x2E50TyseZoz4ZaAq283os9UriEGWU
KO581Fk0V9Nc+UESsRzFKde4StJ4nzqczSPRWorzSczv805tMQf5dSAUZ5jokBo8
cTojRcuMKS5C0oGteGsg++S1oRZT9Kt/e/2zt8/NgE7yvsC293UF5pokp+oHGmLZ
eHOszKp+7syb1QtXhT/zEePnXN+jGBDLSwfRM1dkPo9NUl2EanHpolw7c4QinQJM
6v9WyWsZfpTqFroGRKdCMjKBc3FoJyBU8pv8Tm2oWGp+73V3eqeUpIOKP6PELMSo
xtVF3fndBRxYUaJbKbw5JB2KTz7LooTqDi42baNxK2VFMcFd0pPeN2gCqUVi5pio
amCyeQQYS1CKxrGeRCKg2CRl7qkqpdV47KfPJxdsjb2cr+BOtW+6M1m3dmdeUfvX
mCgOnflVBrCxtKNd89DSote5UilnYsZVHBDF/l9Bz/cYU5vmzMoJS2p4PZKuQGQ4
kPY2dJwZqmHv+2F/I0SARZtFSGj6a5UWO6cGgdtNO2tWGJngqLaCUn8siWKwzTqt
iE7KJK3WuFXti6LaxRe2+ZSdsWIM8GZFuroC2/2ueEcIYkngjkz66/QlMJNq54o8
/KW/2H3+GIrbtb+PtRtVdtgIXmd5/znYxcxV8z3YbP6OlD78w7J5U23Io/8aoWyl
w+nUPm2Jy+dS8pv4tYXirtclL0zLjxtJsj+Ww54w4CGnPZ33YMgpLJm4Qx6KsKQZ
RYLLv4JWMnb6Vc8giU2FnNkH+YEK3q7WGmP8ihyu8QOfrkOQPHi7fQaW2pQAaSoX
+r0ppxD85qWe+dhnIsHkbmnDymfBY09AgoGF8n9XZPH9aYd8+6b70YFIUjzzjrjA
dxWYhB6iijyMrn5v5v3cko6ADAqZpYo3CjE+fki7t3gzWuYXiGiQIClymM7dNlkY
swbCjSmX4mEEKpfok7LNgmmTrgvETYv2rIf0OqqK+Lpaxs+/r0pRk2GR0qsYBSqV
6zE8O6lQKOw6hHXLASeNcyiKUh83dHLkqh2lzUg/pBlC6TSR9vmCBouM81JTWy7l
fe0nLS5GiEhLx0JE8ARYNelnyNGZUsJVUdDkKoGXz0oBYmyQudkwFWuxeO9lP6ad
/4xnNe+a4e+I5spxaMYx3yEXMiM0AgYXnSAa+JEYsTgfQx9n7GyH6tb4O+OJBxoh
tBCCLhPRTqUel2izLX9WAj9DWq33deb8RL0hBvaG2FM9HTMjl5ENsK/gMJ6Q+Ebp
KqpKgQzfWoNtRFB++mSNm6Okjk0b1M9wbfozP0JMolX6cGjtgIXlry31XsWfV+is
PAxwlTmtU16Oew+FOJeDqTmjBDk7jPHx5j1V38HeiUmaget6a27+sVWJHsnW/o5O
JGPTJ2CdfZEl/blMZuFbuMMFdB52IW4j9nvuI5+LNgIOXCJNVwf/u7IWu2hJTK+c
cNLjlENVtVzLrBcL5QFaZaa3odpIPGgVjNr6qx8MONunpzH485hhzXdnUqMgAc4t
UjB5NMtDaLRkyTNtK5J3vmTIBnR96j0ZbNk+/b1gJbLDLXUV3bA+ZdtF9/Vtw1Mz
5kYMQVEMTqkro8y4PWsUEpOoh8It6LB5F1RgNHQjXDEnrevUsELAPBVvpnFCrvaW
iHkIPnl74qZrx8T+dTahFi+4GTl7VofpWiuj9vgwkFLtfV2eSEXrVAN43HeY17Sc
2x9QRIhef7rGmNRySyNnFLj1XZ97btpkrHHFtLAO6X14zuuZ+lxBXLo/fEw/nloP
IzcZWH3VvvU5MNAlHWCIstZB7bbm7AExSAKv6oItN9IzYpZJwLz9azWfZJSl1u1u
glf2Y56B+rMLiI2p8KEEMnOWV/2C4lNdeRI3Zgz7B+RawL6FcjdIE5iNwHzWjV2v
zZELWAtgLSy68uA4c6EBZS2yL3/GFxnfGv+n8Z3Y+Sf5rg1OsEuJ2mAx5vBgSLvC
SY3M45/HJOkaVyImyVPDY0fCVJkZ3Xgy9ix0W6ixqEuVnYDIoyN1AUbxKWpre+BQ
x8gxhZiXnp0aIItNkLzVRb4mvI1AG5C3gHlJa1J0BgPFaOcwEM2US1yVuJuWRJyE
0pJ8DBvfW5iwUbd8K3EG/x1t7bH/Ns2RrxIyaxOX2gS2OtZBhqIkXh7PRHeFT5k9
xY3/PkVWNrMgnF4MfpTLRRN+WtUJk8v0aPE9xYrVznp5seK6m2hadX0f1vF8zU7X
EG+zW0XHIQJR9eu75LyDx8yVKw2Wa5TEBhsOjaQJhZv+HZ75+VDOLcS2lfYZ5g65
KNzcb9q3iQbGLMZ4AdcZDCenQ20HuIngPAK1/XLtt5h1QvJ8+uLxDa7wDXkEAWO8
O9Zdk1SGCcHoaGPN0YYHZaQQ68h/qb2Dun7X/Gb1hU3R/POSnNm98OEsOjBYmSgi
OK18eDQJH4OUdLfZ7Km+9Ks3Dxa6ScrT9fV31FKieFlz7U4DDW30wjr20LmNUvYi
9L72/KJi45xSZYoswXZahB+hSChRlqBjPgDcXMZoN0IcISKSAue51cE55/rA0ErE
LhbrdFHh48OvXIDUw0ylpj9br/TBS37NLJahyDZ+IQ910+/uH6uFcs570Y4x7k57
5eWQC1BM9SWYgdSlJXFtuBwEc3eAoqibrEzcPjuRdydmL/vHThVvV4bts5n77AE3
Q+uR/65SAUgjh7udkVkVtADT/SvdOOZmDGwUS2HnI6nw3pD2DjVrNdUNYfLXKGTC
L15hOXCPoazGMR72kvARO6iftDEEttVmuuHagWeNmscfTnRqX4fTZ2llSL4uC1ee
awiGmYgsvmsXuXQc/HLvdCIvmYDJGsNNM6RR9s4YAgxtmyaMYNV4PwVD62fKl13T
FFVjmdawETOWNoorVYhKpcIHil1gHSi0f8JOZb6FTTkWko+D5vJMm28sEO22yQOJ
BShHx6308a8jMw8oTsmjYknpdISkMm3j4sUKyoLe5x3p3exX2MLeNS4YkeUkYekc
d+ERStXaCOBGfMuqxpEEhc2rXxaXUr+HvNFIW0B4xlMQMx/hGracWElOJ6h9GGkx
lUyufqLXpcoQ0U27Eg9JnwtaHq3A9BwrDL9ORt2Huw+6a9ZczCbRLUlYZflywzAH
iJNc3zeqJHPPm7uXK9xYanmKmYCuUVDFIjmjlc7EAHMWcKjDVxBO8cCnqwvPKid9
c0JDMIGZlimZsznubY+imCrvbdUBbJdwh+kSyhsNtOcUmXtF3u6o5cUu3qa9VpbN
VMYV9bGQqNaxdJWp6aGMSpO5REc595sC2BcRPXRu5Ke3dSKa/LXi/kqZOPakz0Q2
uzCgqdfqPNTZtYNXstn8lU3455Hbt8TuNFP23YCL5JIdBLsZwmsdYFnwhxHMWncA
OoZFZjkiU4sZE783jAIRZuqQ7cBaUTYXJ+rLxQ3IbIztEE9gfRQ1nwo02MilV/cw
NKy9+ATTV2xprGpcgM8lyi0u3Y1S542C6o0zjtTsHIMSGUUxW/FK4xL0qDA7dtK1
F2lETUPyz8SlbnCPr8mia/vM3kG0OFdic2uyTHNqe6svIFw48LT1aEyfa6w1gjrc
MnL/sedp/s0jFCuDFgMn2mvfZ3QK1OwelhdARtRoE58joTvJ+J1xpZqKTJL201zm
CCqoNp0vWcvAcaAKYi9nr4ud5kzEQBoakKvs6TWUxQXH0i1CTHkWyDiejN7P1OlM
rH2bZcQaDaZaz3m/4qjo4KMKtk7+x/mDXqaZaUsXn3TR2nkUWFF8WsSvMHGbwdoo
Gs1r6uXU3cCrKPEpZ4kMRwCn0A6IUmZFyAgK0GQG1n7ifGkkfttmvjKt4yM6mL8h
uXE7dbxC8jJy+U2jNCKnJ9RD2EvRO0gjpVFV9+v3n5FBHFGZIGkuHDywzsDRaoFx
j87kRIls6KYH8eKvEwHvL6hKC0ujsCQsYwx01U3HLfCBorByfLkc0ac38QzGjdcT
ojm8ibvUJa42C72mo4EOU6Vx6WPXGfCXSUceRx9+UyArzwLdm2gWvvKgSlcq9Vc7
Lu56mEotvrnZ4R7ZDW1SLWh+JZA5Oxk21Rkro2VXKzzLRK/2D4alRDr8wL4Ldptc
r9EfjyPr0Xl/3AyVKIPkIGwvIsD/tUGH+M8TaXapW1e33SxYCBimQ0wSDDWsdWUx
0dYii60IDvv6H5P8H3xsyDyQw4K4mLJShGVrAbMWLxyZUf1K8iOLd+0eTYLm04lF
nyzo6/lbO2LSs7f6hiRrukqq2JoROjiLMxQMbDP8vZaL5YLV9smezVPU1YG669mK
asD9k1MvEp0nnJ8Eg9icHJoghFzwx0GuMhpJ32poprMpEKwFfVCwCdlWCsljkA6R
UCC/0oULNpPXHlhsxkTV2G3X9EDr3usA7h5L/O1N+n0C30UYudBhUa84VA2E/lXh
dojqtCEAyumMf1R5881LCfFqEZYuMQXV4W7dWyhZL9wsBV+Y/LW4KNL70XltzVPI
Ypz2P8n1FGFpZzBzd7ZR4xbS+FtsUy07lBRc6BhP6yljOBmNy8aF5orOIBD/OK1C
0tAkEPJ+h4SIHXkOXPakQyN56PnVY75NiRnYjLO11XP28k86k0ZlFl82Jod6vcas
FhSYATT4/2ml+kJhTdOL7hNDRjBLNNCTO1AiMq/V6RS+pQad8SyGhhhCl2ZoUJbN
QNg6H3Kf7lSvKjtPNPtAAzwqi0BPyUJ7BMvanqbWrEpGW/Rv+nOR0rQlVD+P29Q+
dYs5y9QZHaoWB0H/LpMa4C/X4ub+or5+M2SYeJdrgKaG1X0XC30NDktS1vt8i1cJ
xkD+hG7l1Qj1AQSeBJ/HzZ3LNHY7v2av+81p04xoKA3UZBGmncdWphCJwaGkOQQy
h8d+CliNPblpQytt+KkSKvajrkkBBp2l7oEzl42gyaff3Hb5UlWZ9eANeRIRf0Lt
N28YTrat0VVcHjTfIfyTgjFIc9AmHy0ta/bsfW+kXnx8Hn6FFvhP5ioPG/4M+vJZ
pgglzDYjbGlxfduoKM9ciGs/USEntZDoRRno5WfoeivNcTPcXx5olTVUvN9A5xuC
dJTZTzukmpNo4hxoAUNo1VEYoIen8aadXnL7wSHT+FNBOdY3WswGri5YFr2B1zx8
pN+MV335pPfRs3Z2B5BUDcUuv9aS2mmseK98aB8/Yh8TlaiXq9VK2q24O1xYiIeV
+NmhLWwh19Miy6S+3Sbulics7aMl967efWLA4qSGD51Ofp01N5+gkqZV0krIrBcL
SjbT3LQOJbkn5YTYsFbhmgyB0fVJuKzk+lM9cvZYfeUks60o9mhVIEP0xghKx0dU
8ebAKx88tjnPU3jShP9n1TLHsP7dpC2ZIKYMnifG78433zqVvgdLxMRGrjbdwnO2
k4d5b9JbVoqGR1hhMWoYXPVKswb8ig3wU6HmATvDZpiR4ZFLtk8ahgZz8xBdikDn
HH9Vq3hOf+9Scg04foa/kRzaUWlM3tMCN+kjExIBEJ3BZgzskAswp8RTouBgEf6L
Y96Ll1ml9Ghqa9T8OJlw3hymqLd/b/ylv3bWi4OolXBM5FhMAUZyTU91N2LQ4rGb
D1mjY5WYHKQcEeQLL/B7AqYSgzDMdGidcBxlO1sRnfucHlUdbjD/E2BvHRQAc365
qr7xgdiEr5gnSOboRseQeZqUYWTUwOvzRBEwoB2V3VwZqgU14eBPh+l7kRUu6fp6
EUeKbvBgVxX9A9E3mjLHqLtuhc2Fg2oR3B/E+gQUmgYT1O+vvfSb/lbio20fy+tC
dRYbBW1cUPceaY0ImGVa8LqzoQLmO8RbmHtxhIdxlHOEgSd8Mue3yMlITLLUS4ZP
w1dyPTcvn/Z0PS80KelQFcKnfJ8gccaTUhcJ36+b6CRWqAwpjYAZhGlOzuU60Df7
v1UWKllnese37/kxkJfNuc1yagg1g07Q/GzOsuyrHuKf7uVflhBhBy/ScTcepKCk
oWUCLPGrnhAIwVBPIMjptIdQyXVT1IMkogyIilOvtkiKtEZzm0KKqSrLb8XRK/2D
NZvavHZHh2x0ZS1gw4PfQdOttpR/SJYeZfcwunnhFMkuG23NT/R9Ona/Sdt7OySt
AeUJKG9JNtOud6479+pujKQck7hkpo1LLgz4zjfzIsGwtNDNAcETBC6Hh66LHHY2
QNstbo6rbRAUdlrVXUsxc2nUxEy+jK++9MQtobOthm2CZr+wq1a13WnRcn4aVxG0
NcmIKHoLO+L7PORYQygKydVTgMzMoMFtTUYGyTs2VkVQfuDPihuwbOy2PbPi6i4S
p9znIMJvMs5KGGg+6qwytkOV913JiCIQcd2oBQCk1GoRqeT50d3cY8/+VC86vzRz
yUbeQ/Of+yStPoVMvdEBv7gCjc1QKcDQKBUodgPqYkvTYmKpAy4WoMb6D4V/WjzU
d/NyhXff0Pp1vqrazg/9hUV8/9j352YkzpIdgCEYgmr7U520YT5JRLf2GeWXqArU
HJ+UQqyzaWShdc64CfjaHYsmBBwPnzWPpcWnXeNOIBT8LcA6FXAVGFy/bx1mfV9K
eMJSwuWT00M8zE8fLsq6hitxN6kbG2b5h1JiI0PP4B127pLGbdUCtvD87m0XHEh7
0m6JXNDl40dS6bZBXWdVSMPzPKZ+pBX/OXVSa6/REfisUvoEXMlX8ABbuqEKzR5B
2eGy6aeFGt6xojGlOkB4fmNCug33LNLGyliAKnvKzaVFOTvgxSt5YvrLcgOeRLBi
LezQ3F13Mhehbi+AyH+NHE2c7cDRLTR1lcz69QUN8/KBfqLUmwOi8Usq9qlm7KLZ
jkc6L+y5uHhPCA8lq2pnemDLdtd260Ob8TMzTKlwmXO0xekM4Ws4B7S2JEX73W1L
9DTpBz7R6kPS6NzN6yghhe7oLrHB8yO6DaYu6mLfHy04EiLd5/GWWOi3DBn07zyl
EXhHZDoJro2pua9ND50FSmtKmAvatl0+nQSwoKHI/EptVkScIjENIxfifoOTAU6/
ZuPVtjM18DGSkERDszeEpqJBZv9Bq3vMosPufuyHuNpK12ZCsCKLS6w9I2TQABY2
wJFE2i0ig85E5ERLT3GyNq0FDU0zGNhIKZzK1szBBLxzWUkZkb6Vc/tknsY9PSyD
g0Y/mEUro2mIiXdacIwQWQKTuY3gB8HNxpcpZV5LvuztLg2fcNDmb6WdQgGmWFcV
hxngJlGN5hyYn+nAI+doJYQ22s5JznfaF0ZG+SFQDZUgBKpBuQlRMoThsuQTnUqL
d86WZ7JQMpELowwwHGh7xBXIYRLTvnlikSVl0e9MoE8ZhFVbgjLf5sEp89r8BaRF
yfChGQM580fIer0UQ0GXsD44dDxEtxRByAu4bD0MI8ggllylwWDoly9lBBRjtp1h
iS9K9uF+b9Pl6o5sBbUbdtwuO96unKEkMGHtNGS0Bu4wFYVirqpp/QGxzB5Wg2c3
1PWgrJN/ZtrDTEJ3ODD9cvpN4PTkF89NjNgombPPFlv87oLoS3jN3A8E6t3iBI8n
RcE858UT9IdA5GZwdfu/jq4uN6BOQWnqCuDhvW8NkGJ1xX1/LtIZKxJakiGwmz1l
OEEp0E0KMzHvAsedMCLZXSKyKxvvouRGfsL6ecuUjVjaX5fH1rfhv9oY/OaH0sWV
N/23TMh+/mHm+ESf1VKOARp3cDAYBeZmCjU1+sghNFmD18jIkp4laws9k5Z8XUM3
4u8hNapc+6YqmtUvRvAUfgTbbXoyyy6CUU//wwsQYRazNS0e6bTsZ6I7SZ3q14NI
StTVaUvLM/LKaiqPHPL1cxFcBMBNcF87XKel7X7OsVhKlG008T6EQAfzBSXX9qij
ZSE9qSlF/ir97kfg1Hk/Qe2O2Lt5PDn9CAFJAJwCM6VOvatvCcgZjwU0N/a8fXZB
q0D2eWYTPgLt3OnhzaglPQSQY8+nICzBta+3HDcrVTzPEDqpn7VQghE4IbP+YzOF
nU5MGJMuJSs+7VR/m+K7u1SEM8OSvSlReZeJTjazmrS/5buO2joof+OVnygtvpsc
AM8IdhJJEoSXuAff8mCcAvcVbzbFfDMbZdXiKqX0SO1c//imIaEwPFlI5Z2egNTF
RVMIG0eGi13fGAbMC0HBnEfnBmzKpxHuiRwGswrgwCQhKNou5KzteeqYENhMkkJ9
qxBPRBY3XybLQKqDDIceS1mOOXjLLeTn8UEc8DXK6mN2AwUvS5STRGmoyNGNLiu7
aH+yluIxaJE+r5vbjJm7cI2FrIKVOgAEjExzG32BIQe5Gwnbt56uLwCMhPvvIzoV
6SLjrVnLVO1dJ4GazJHe0Jm9sDIYDKAu78ylC4773n+YtTFQYsmHA7QlQTqDotxZ
/GHySC3c46L4ku3r6HudsbnLAAQd4bf6HXXNxcM5xeOTmoUPiidocBLU9e+Kfk85
W5pkSLs5fSe5wMQ2E3xpCRKJJxQdzMPVBjTJN9EGkPxxo/KAp6Fa3klT49ZXoMGN
EJWxWap6aQ1bRI+t8SAMf2XBu9XJpJpCLz7X8rvZ3IMWiw+WybkDH2ELY4UeuMoe
VDckMVHID2IXCjWc4Q8fnMJytXW/LV6toKIjlpn4+VyeHu8F1DGvO5QHzLOpl+so
3evBuRUyfNWalBRfVVH8eFP3uYgCco0SKu/VXLfHBwDLLyGTNLBsRLbrGdHSurGd
YKKxt4hEAsFyuvtW/07C4PsmCxMG1d6y2d556h9HIp0nxLEM4fYtnr/zHsIpWWOQ
2nTs8+vdTxkQbzrKmXQFpnpX2n4P2zC7rpmqf1z5HHuEfAhWpxBgJuupFLgljSPK
lVm2bn6Osm40Gr5fnS3sPzbkT7Xlriuxs5rA55Id5FlYq6+ToJmuMW6mb0qR8Vx5
6kuvyZrzvr2OeMzNddLC7u0pQ2zNZh9z6fp5WBxtMD/WaM3rhBP2EJOX/DVSNKF9
gGT8oYWqEteObwIhN5GZ/7FlHLr+V36TBwl09v8ajfH20uzx/98OPsflOmL4FaNQ
S02iq1tRVJlfq6JaDdCuRKrPCQpwC/LfTcPNi4dy5yareJ5oXfBlYtZ/sJidR+s2
IChhbuQFY2LOaDy/4tJ3OTXFmcQTNncahEOP32swnBtawr/Sa9Qvq48Q/zzBhDEr
AJBqzfRo4SRuk/LaFNbkEQHzt003s8m0yPR8Mczq5crKZAQdkMAx+Cw90j3SLskO
1rDMDEoerhA8z9RVN6hf3JlswXcN5Gx0p5N3VJ4iwB0zW/etTfmsnqU63CVGZJDE
FYf+lv3Q++eYzTHGA4rl2fyMiAGvUIt+i9JWZG6i552DRzypZmJaaPLo2rEJvKuh
iQqYjkBzOFYTNuYWs+BcQGFiglcpJ2LTNMOGdEqRwGnzz/YUKpQOsq5m0h4VKOhD
Ub97EOUVu1JBPeo+zoGHtip2FfRMeB0Nd/Orss0l28bCf6NxQc+kq06Zkyem6GOm
vvt9hoMy9UmocLwfUiTav8iLEhyczom6B3ISgnIamE375715dMD0h5EGmtoiMNiQ
TjKv3Dd9yTYW4sWQCoBO6ikb/SDhSLL5dnkcTtQ8I5QKStcHMB2LcEbPxhok4LND
6+aIqS2XvllZ2laK6t8JJ31hhAeIX5o59MwRy299Zi7ZoOzAxr+IR3NILOwnqmPR
fDxZi0w/yZHT49PTEiJqlF+WfW/5poxU/TC2gmqsKHd069OV2DE2aKZ0+rXtipeG
a8SWgz+qKknbUh0AdWXPNhU4P5qxHWGSYdApX+48L0Mzzi7zYPzhJ6VB3np3bB8s
yhrWN4atH/rroxaAj9MSrobrrMnvE/L2Agr5548ZUyLohjzX4z07D3ReW6D8XZi/
NdbT9uX1fas7yKkMykxpUB8eh/Qnmgs3UdeKVYTmZr74FuUxGqvekoaWTcEgOcRf
/TcY6MkfeJnXjtDQ2YaAFpS3HS2qbq3I4Y1bphLWbgUTbtwqr16l8nxo/HkLa9Y0
mStHynlYXKwCWWCwPqzx8NsSS7Cnf/lXcCCP60q5oyGas5pjkS1H5GnzY8C2Fs0b
oTEvlbHxXQTvI6FqeFL5li7Apmgt/vY4cnY5fx9IbeGEVQe2v92HE+XgcfZZe8Zv
IqWwLK+9hBO9mMKuSd40HquAyORb1me04O4l86iywpQi7YEbH//aEJARXlTqi3lC
6zLNiIJwJSSmBN393sG8kDG/IXBzeCePyx90L9XWL6wAK84b+w97lwAVBu4zgcB/
jYB+HsgNAoBAuwGcsAsmd7on/pk5ZahedFGh/X/KmTCEJp/QFlCOBY29J0GTrdwD
pqAQhZdWDBPg0tLhk3lT4wC9m35EXMzQesMUWhsflJk6tjdTZuuEoZ5KMcyaxRnl
LGcofJHEjjMyqPx+nwdJbEjQYOr0RcW/8oKnomgpMa0YKCM3LH/+iOAi77WArIP1
cwbRwr1NkBT45gjHmtTSIZLzpT16yqfh1yLDSvtUv82FB0kHXwNuLnq83HUOV72N
HY5b8AHlssM6Y5RworOMuRy/TiOAAmLKtV14hKDqKIKHS8n6BgRgflamjbGMjcRG
dy+sPY8gIN9DYm14liPdKk5jZjusA4ps+77DU2eflJQLDd4LoTwOMfc0+TgGfnsV
sAL9cMrJms6Mq58XZdg+r0/QrMJpo7HIw0ZhCzzMKzLHM16WRIyNLSug46T6a0Qz
jXLwuK2fnyz4tsXZudQfievNBkWTqlCNAIfCqHZ6VE9pfK8CUKuhUd8NGZJzR8RL
JlTkziVNkaKOqm8gOi6yovzw6PJrSpRmS8ZdUftX570li66t/OYoqpAbfAqEn0x+
NibQTDMQ0/KPtriHKkoBe0cYqEgslBphnzv+96xnVOc7nJiEBBQs8fMFkr63osqO
4lYBVgGioO0Rdb0fxfUmzXUMvmf3JVwZ92SSG7EF9MH+LdVb0n5h3L3vC4Cfe8BB
kFoBq/HXBd+HjZbTVJCLJEthtHSm4tt4Ky+cjWsdC60qJ7D2nGrNLkvi79zCIY36
7L7XDjHe4vNwMoN+HWACE9kZPblR+n6i92yYWqYmSZlS8WjhXaFNi44k+cg83cuV
9lD3bEjdtso/+9t7Mz+rOSbmbFxxfP4bLeoUN+4FJDMrNG78Nl0wNAsHAZtRtzOf
E0trHC6HojZ1X9m9ZMQOSqZV//rxK0B8TXeeGfhvok7VMqnE99Ty2vqLpyU1Rb4m
b0hPnw9jO4quhv4FYLJtvEX9FEwsTBPJMR+wY5Y9eOSwDjnWgHIVym6ulM6Xn31r
NDE7XSKshLgu7dRdq2szB6KVVCKNOmZ/Aw4pxRdUf202ogr1b/rp7l3P82bCQ1za
7NeljGC/jQWv4A+HFHl8sEssBKcJWdrIZWrzWKH1v6DA75Q4KTblsVfL0XsiFajN
Xj86XKVEUba9POaLojxFycn5s9HFf3i4AcuGGsXFTEQZx8vJgDGIk6skYGu2CqVF
QHzw0SqRpx/ReAhdnF6w0Q7FmCXw3LyAJ+hW9L/y1n5nBgw95J1s8n/EscD2pBCt
SduSUvQbIWmXzRsytO55XU61Zrk4dyttS65f9lU/jr4soXP9dkgC4e4lMp7o+L4Y
VIUUFoBMhqrDxeK6X2n9Rp/wL/rP33WWHwhvnEPcvoq03hR6Mt3+RekBwnN1fCJM
w9DYf6jm1+jVYjg7TE5TO3y5kxOfBYl0cwYcclHBwaPMi4X7HFFI06KawNeJVuIV
uQA4XbIBj8wtyl4+Z8sQht41TyBlG8Gvj+pMxPFRU82oNjW2IBdtepHVbrP3iReR
CS2GgC40yEAWZVAwv/xo+aEqp7JBxITvAPHGyAuFIrB5+R3JfMvyH9QuUKUlfYQd
USf4gens4gzJ76lh68k2l/EuxYDt2FvE/GK/TPqHFWxlGE/Vg76FY0z/428KSbxF
vFfQaBEANiwE57V9EE9UKaKdpgqbYJvfNT/RYYAu9k9815aNa1ZnfIVVal2YZUyW
sTveTOfbuwIuDTVG92jcypZLbbwoZOq7ncIvNEQqCiEWOS+Q2SqekgGFJH/5MHp+
QtqZHhZo//dHTVDmuLE/IA/RwgCLNssNWw24QZMxa4MpSfBPnxlHWzNaeFpcCULw
GN4OP232gLsO+4UFQvzF9SjHKQLT6OqKfurD1fevJDpdHiKfI9cIaxRwDC60hQEr
RVwZ2bVf3SaQB7YDB8OuVuDjsPMUeukeRORq1TaDnI8Si14ks4cMwWiKcmoJMfaz
R/w8h3LeRUUu9ht0p1NGisGxS+6/MEHJyFKVkvrN4Gfuwpg16HITBOLGwjbH5O9t
qDCn/5emc7cSkWqsxSJkH09g6T40a5q0AnglSB3rvViW0FwznaEgiK2DCOFJqrLp
0DL5/8XBsbOEevluFUJ4pDEoE5b6qH1Ay+yjp4vCaO+pVxas+ov6uko+8K2YaKQZ
dnUuScpN5+SRs2kCR/qsCmip4LCd962U4wdem50uEDqRjQnflelixTiupoFt69WI
/dfPxWDEZcOwTmqh+z6mFWgVl5eYYab6/tZTOYUlyCMdmuL1Xj/jVK4zWV92qryi
UcqJuRAOKEnmdRZsfaVhfJVIOyajVNMXuJpXwBzBR9r6jK4e/M03nYsNCisw/hii
07ZMXxl7Qy3dvtpc4s7f96p98baXXqpsbSOnXxcLyMki/+veiUCmyr2cpN5Gs+sq
pl3VRy8u39ygO/FxYESZa3i5RrkP6tm7tMs1W1LWFxsnkyTehXZoe5a2AJcfm3d+
aB7qmRdbxfhDcmb88fO1dD6dwO/lvfDh8cih4QD/p+MbMxa8wA4pGR0LJCup6tBo
YFZrt41gfYCMynK8WYIosEt93h5Ypc2U70nyv9mkfaFBKuTiJSaPbOHc7g4hJMoK
YUio5kTU0jsWnL5ok6xEJXH9WYSzIu4lX8kdhiMt9s25di61rU+m9vxU0sJN4Drj
eVO0q2IfnU3pu7SJ5+20Iy6EJoKmJYlRbi/3iE0Ajy7DCldFuNP76EZdvPz3aKcm
8lU+a/9p8LKkYxtAt+a81BmvtZ42czENnDsaLgN01iFhGOhxtocM80zW83d+ujm0
RprULtw+0W8gWNWeA/Xd2GQUy+XODd4LiiGu7M51Cxj6rZfnJyeKyFKQAEitqwc4
bVGKdi9Jg/LNU31ntnL+WU5Pbx/EA2OHNzkjAf1AYjXldPJ+2qKvVl31iBjflA1O
ibjO9AR7b/t6pwT3wgH8bA38eHyc9xCx07gZ6aXpHHEWBzkj+whzstscfPIDejsx
Yc7QlyouEq+8esbzm5IRk8Dx6g/j2Ha29W0/mak6Gvs0FxrmZUsR1bTXAfS6bTHp
4fyWIX3mzJSKgy8t6fZI1Dj+EzCOCwLSXUZGs0Y6T114jXjjN3KMfVlpty44vtG2
63SdJPmVhKEnuBlTVWn6pqEpLhG8YDsThs0EYr/HRzTtJmHcOik3P3aM/xB2L+Wr
wTLwtQsjRRosN+brsnC82KfzkyPfBsalU9vyZAb79VAIvi7zWCwL4E44dyG3D1IF
Ay7NRu8fxdcL+a/M+2u1rQ+xiZwtQDc/rg9aTyC1ftZkdILxXsRT9mnRDkbvu+y8
9TKV5bqG4cTLokzYhEtBDaGP3aotNg+C1JQTStmqGGNUm3QMkRBb4MwpJCiqoqqb
iL5DuKJer5KaSIPrTD/V55G0vZWsbz8Qr3yXIGW0AnSjrPAvqQ83CPLFhvEbm+Gu
0MZs07J39dX2ZOWgXQEj/V/u1vJ385GkXFQS8YZ0lG2WPJoRIs3gi8klDv6iR0Z6
hHTuYGfm4l5ZWEAwAkLXLyKOeQ32kTlO0Egcwnqqp+hyq+fakjzZWd2IbTfL7tpr
KK+tXOHiuueaMA+Jk4jI9Y6Pz/q0aQu3jb8kOInCoWm7iRcmnBm6Qk1noKlFtmjN
zwrx64EikQcp3WxQLepO+fM/fdusaWihBtch0pd/4pUJEGRUIfgfftxfhof/znGO
OxOTf+GezpsD+iUOrLIvONLpcMXkpfkIX07z7ctQyBUXkfItALH6HJkAlSLlb9iA
9TWP4T1hLLNnkrRmUBNHH4mxMRZiVa7hFhV7xPE+Oj7ryGBJspJ9uDP0LMIvRjMQ
m4vXv5oyLpz5MAlu/21+/74O/TQ62M7NqhVBwW1L/ighcjTUuflRkv0KEwVbCWtL
Oz4eEEJXLje/IAXe/zdXRjnauhycUXSbU28QLwOgauytYqxBOU9D4i6PlyPUzPGk
K0gi0dRmK4QGhRrMqpOir70M170rB54PW/BrFlWjSB/qcWHZDDFbTeXNgnvy97Y3
6K3gZ3WRFRwbBkmuXqe/xSjoG8GfTqaE5I4tGF+CJkXLAeP8mxVT/L8dTB+Fi2jI
rljRbOEOrCtu3F6irdG1Q5WisVEVchS7oFVubxvG+nAJFSK1gPEKIn89KgrzRr/s
z4eMxSuqhDFb9T22TxqNLeK0rk14FsL51HivW7xWHUYrKbAB23FyI0GdWg4+GuOb
wa3xj11CP9+g0ZBMmZu3GOfQUK0zeiidRC8RshE0Ign+AeHuE0lUWJMFMLU4Rtjs
RMD7/YiFfSwDSow0f+2hwR4iQIyF17iKP5fMzYJRbPj7Dm5q/J3H1dxliAch88sy
IB0gJlA1Vqevq07MwJjVRG7uht21OaASMmypVOyTPvMkDyQ+XXLtEGNH/+wDXD1+
AsL6TUow5bLts9+vu+LDaNkJGBuevx+A2oITqci4uYxULTlGLhdREwN9yg2RYpSN
qatxOF+SRF1UjzCkFMmwH8xkKkD2l7wHu8DBGb+3nSk4ILhKH5WpOPl75bDFXrSL
2nyKiI9Zyk+L3uFPA3+7/lGvpgez9U4y18QfH08P8SnkhMYhXbyAg2deQCf6liJf
ego+b1hDF70c7hTuwcDNfazHNK/oRvvXCWHas0eQQnOZ9yUD/Pl6MtY4PThu3h6o
JguSPMFIf7WVIeqNQ9PlLKkw8+6aVIYxNHFH3ysHo46yjkv5lVfv0ufBg5YryOp5
/wGuiJaet0m7wpN/DrTprMWR+nKQGARUpTZALsQ4Sk6mtDyNWhCV3wFc0Z6ufGFX
8GWGKMnG7DAPaPOR1VgCGLB7G4Qhx9ci07l/kIcRXKHpS4Emc1UQUZESF1I8rfvk
tfiMKOioGEmFj/EcZgc0CwMBPA0GnI7Def2Y4aKCTNA7U02fBYIjkUdt1OYCzRfe
3a9Qptt4LftFkb7RNa3zCehOJjr1Rr9IeXQwqai+g7USE1wzmPW5D/b4AMm50jxo
316/lnwMB5T2MFmMKJ2uajBi2TrH1/mkRSEBwD9jXl9F1dLnWKPZP0RPU6g5o+q5
sSNa2yMKrtt3HNKn+Vyan52+UU1hzXZBRNXDdYF4puZpH1+hvr7Cu7HzcYTa10N+
2Vu3TFm1jHnK5+Yz7i/XTv99P+1WLISRe9JvXNVvtzcqI8LZRKUtJhaWUR38OClJ
/jKhcyq+aAKaIlRZDVX8fXbs2ErVm+7o5hV6dtQcvmY7nykFSuaUCuTuo7t2InL/
nw/V47vUyQc2hENK2M4Dab2DQeQZPmCVoF7Q2xO6ikQnTh9F/8/iCFl5n9JlUcxK
HJ+jUV46gBdtW6wdLTSlRvEaCb+/P5fz0q9xxfwf2nzwV+2J7YNr1/rpnAjCVzCx
Xc+Qya2gYeRKkUvdWsaS4vYaDEWyvwFhbhfk5BQ8kUBRls8NF+PEgo2zP2dJklO7
0vD3Y5Fe01rrvgpt9IudZZgpBM+Tbpe57xLaoOO+LND5KwZPTRgxFNhlqkP8SzyL
f/vCSkn6kMmGKl2hBBfL9IhSDDTVYbL0PJqjebA2oX0qLfRV17Fdi9iE9BcjFkGm
vC5ZIC70R2zUt86ikXnX8cqvTqG95RCZeKMgnOgWIOGG5LvdIDD1kgCakUPsG/Ul
61gN/CIUcFr4fbUMd4Ys5tR4ARwWBEI6HKdfcUXdyL5bYHUwaESpoHB/UVTckvqC
e5TPnBb1Bjfex6GBw1Euvjn1rLYmo0cONYRywBtiVLONcJxrwWJL9WmqOhC3QboK
eeGFEem4C0+uyCE+0elOJTKmYQqNlv7/fNWnf0rDfD0z/T6AgaZK2zSb6KONY78Y
uEFrTr4636H5brEqBOquXgWqcK4ejKDLhC6iwzSmST6RCG4XicPkkkT3pLVwxVOY
cX9PfqGMQd5pa+r6CLl8Hm9rb0plH3zY8wrxNe4wEQM1spdCSllgTlp5sGDs8gIj
t1yuuoMf3X2k6xRoKGilavLsZEP2AKBBIU1P47lQ64c/JwD1KfA7+hygzhkwGUZ2
AF8o57AbaqzusnfekbdorfIzlRa6R/AB3r4NLt2EQMbvjakxX+68n49p94mt5ojF
2lg86iTfAew4AbULkab7O/xarG5FUdmwHqB3qu4DalZS9pQVWLHlYhV0z+/Ib8/g
VRlQxoS7run3a44EhX6XqO47KjT6k4D+MlGASyQEOf/nrsMCY4K68e33X7kC2P0r
EvXZno6dJzQvaubH6qbPtAVqh4ZdUQuJ1PkKOQ584QtQq+0Eem9BZLLI6X6WjXTb
L2eco3an3Fm8j53x/T3oiwN5sml5zIy1KQCVBE1bhjdPFeOvlW93crWqoAhxk2bv
aXpqKOwP02uXdwpWi5q2Y86OObL9T+L+kvX8/6kqgNUF92kgavJOKB1IgqUilBzZ
sFMHlK/IkWzBpJ6lITpxt9jVSXUBDRmwPDNQ6bKsNLDAN3rxzPRK4vV0m1obctYi
hfJTr9UOwNZi/1nQsuq7u4fKaouPCpTWVozgpBmPOBy2wxub2l8tT1CwQ3+3zp7w
m8KRugUFbR670ne0EJpPeNmjIW1FWVswW1yIAwdvpip2G03FYBUIEhxJp0zVZxgb
M08pv0vnDxWtwVA+zSAz7omwJ/QkDT51JMXl/AgM8RGV9irPS7RKMLe+Q/zpU53c
/XIPaSeCf7DiRhTantuneeebIUgg0YbHvS/vwJzMe+0PlANX+N8ScekhtTWK6AFl
GAN76cTfKIY1QWW0FcumOVyhtGb2v74vev9r5LOQyWDfwfnG68qq/0dWvrg+l5Xc
Co2QDbrK2hOHnWiSfwd8JkeAZSRGT5VoPyiRxNkYORw4ES7pG0phAqYlMbN8n7xc
sENAoZWURinqquLLotbQ5QpvdZSh7Zz8T+cDXw/6h98mXGAh4oaiy57oFUTAbhwg
To9Uxz/0O56+48HrN9vCr/STRpZH0g9JUUO+RbKClwD1sUPUgpi5ASlYb/y8CboN
w9rk5Bp3NvAqm+J0QS0QVIh3cYP3sf1ePzDJNqkbdKjgXjzuCO6K8tacCc1IaFKV
4f15S/qYqbN2qG6uLAo7MSwZvBO7OElpAITep02MjBR8Q9UOQo9yOfDmQOjjXv07
jLJG38jPpUETdXPsaW1XqDmbDu3Tqm5dMAdk1MoQ8Zxodb3y3y6jDw3Gx6mDuIMy
FRmRK8Suqbpu0GPld2k9K4XZKcFCnFY9kwt6RNFJ4srF6sz5oTlCt8FSSAOYxXkZ
mYVO2aOuI018urJ7u74V15Q7WXXcuCgArlX5jgfCnncYzWELBdn8MrZK6+O4XHIu
EMehVHNBFEULVc1OnlOMdJqj6Br+bu+iPrF9gYChVp5rPxrF3cvvsDBqcH3o0rH+
C6iRSBcdMeXx9l2iCVgbUkqZFEcBEXL6hoV8BLcFPCYO0iBbzR9ZK6ecgZ42aMsc
3gn4unzLtvTSNfIxGDPQl2ZktRl4+Dl9CLdtTHIZtYFuCTpFF6WxckHu+rQmC3Pn
+DnHocMZKf+RgN3b3M3B50MWFNFmf4xMBLLUwvtDeWs2+G7BnWHpRH9uyS2g6f+u
c3l4iZD3uEOFp7doa8bLl9GJyRxBviRGZxvuR4L50HDIX6SVYN4LF37W15/Ix9qu
Hq8i3oS5RVe0SQd8l8QjuAeTQh97UhvOWlwn1K+QpqNTG1NOBQ1IviSSr5+4uAXJ
5fDaMb27ArytwmQulIED746FQiD+fgYNCja/psl7F3rr0SvNNyePNa3cprF4FbB8
y8XnSQgyX1SXIAwo69iLlVWeMzl3ccVVwJ2eBjrddhTZn0EMaPO62z+EZ3WCCIGa
i3Hfd5nPF9C0AfFMnZQemQZJCbr4To6f6zZVJcpOdPfp50AM+qlkE/5A+HQpWKSR
mzkFL2IxSFkqyeR2GtMWCzlTZY2sW56e927IIfL3iiE5uc3VtROYDmneUaO8L3IB
VYbk3AxGWqe+ARAh3YGb/Y6i0AYtilIyszKMURZeelfbrAootmwzNwhd3HykaYo3
dIJnMHFxhvnhogwzCOZfhokRHkge3umZSeB0tauRS1Hs6lAzntzdQDS8KHcSCkg4
P+rMPZPSLvXXgeG1PV/pH4Fj6PrO5rHuAbaiOBx++If75t6OmfJaQNhka30Vv03L
AEa5Gar7TcO9FaD5gUVmgaBC4dUDxjDbD+CmZU/ZrDNT+RcC/CzwIY0Uq0KmrpIm
HZTjkHHfu3lUhA6lhEJez1pU+atMGm4E3DmJ+S4gx36uHVdrN8kgdxc1HFRWHJC/
MMA1OsxN1a1bIF4LKql2928si5qrvAqHiPl1YHlc1fZtoezQp4kHZDcPbSxtIwYN
JE5ZCfjWma+OsYR1+R+ledvSHW0+U3Y5Vl+l/Hy1G3lztOKzeRlmvWT1Xaqa6GeM
ocSO2gv3qwDcgh2tcXuHV1SK5rLxbV1HHMaKljzE5wJs3nS/xquKZZXqd7JQGtI6
t5LtHPK3L68J23lRv7n2JQtGeF1Bkk6i5Ao/BF1w65kl1hk+iUwUARZMJtPb3Eod
VS0Xly0TLdVX++0xDsL0n2YkSRN7tePbKY6ZDjwPgPs+vZlYAiH+vUaUSwZNudJQ
1Ln7joxrZK4jPtJKoPFh83EmVQtXeVSEctIOEONGnkZG6zhcjFERNzIV8icp8Ji/
djyhMU/p47uTAAli81QBOQEN4X4m3uvOh4B8q9B4UH5AOumy77OKrcXSv00d+oko
EGL3d+Ak3hZQoI/BOpoTEdYqv/ojveujYt964D9hBIsBiTmnpxZdc5Fhwhh5fdHe
dYS1YDD4nHd8ReTPwmYfhqllQHIkalO7bAqQBh02Uw0n+F9uCgi1rI9kwzMEbSQJ
RVn9WZvVaZ6124D4JMygm1wyxPEQbmQZpRzHOi6MlS35RRjejalG1aIa213qyc/P
r6jl7T1RHqwcoypTv/J3MGB1OWrnhCHjyw32xK3/1zlNdgam0F4/zdKNYptwPB+L
SVEjRoaFK8D5LNHQ3F3mQ4Hyg+VE7JEXWSJHjVZcW5lTuhQZuKe4MMJsfm/LfZoE
fKTf5SbAccq3VRjSrHK8vScngPFHKAGI2be8oFKwF9UDVabBSSUhSYtByN+NdieF
igTGcb8+sIVrnCE5e6KhYTUMRu5N9XwYWhgHWeDdx7/Rr3/ApCJIrAdz9FiE0jsK
3zmX2ZUJ+vuzfWHWnrKg0is9gYYIYN1bl39uks/mCJsLu4aVy0PITnTx33T8S6Ux
eWVC6MO4lm40LvZHkr+5PPXomu9RBNTxemHLSGEXGlnD6Fy5vmsaG6PJZMH9DE3l
SjAGn76hE7tifh7OWEzFOATsWiH8dPhVIeP0aFNvfx6n/Fx1nSpVl4hCnv6os6Eo
G+iebid3UQRFayfYvcjZBSof8Zg872gCihn+TWrur9E4a1rjqvw2nBnGF0VZzapK
oTfvavGaIWw3YcY03WpOA2gxtdyQuwZj7uO8uv5JRijj4LpfVbgeHfdAf49Stqg9
r5WxydCaeBDMQ6Q8xBDpTS0APiRQponPo7VofESZFsFrnVxogjQzdVnnmmFllShZ
3acm46tLGdCBGx2W9z9gs7Hq+4PMLal8fMPqefhQPR0QvKf3TNH5odcD7Ms373H6
2xSRscnk1RkSjqEzz84hvUByg8kjXLtJdNdbzJY9ztXQ9DBa5S2lQLeOPJ9s+BOe
1Wz8fFLPX5n5Sqn2vbwTEACoiq7Z7ciGsfysqXKGCYajX8RbMurTTeakeOeOM4xP
Ra7+kd9IO25PDoJtYMPRGg1/aoqa7h2CahQPSgWAwDdDBybN71CNEnYK+d3kwEEN
/T0RS+RwxbacIWfseJBXzJ91f4gmnB26RWT8w7V6wVOfnGY3ny/S0tl8xW0LhlTA
n3emddTw62K0T5trqHviIsqM3Ma8F9UlEOWq08UTNjYy/QsEAzWHy5qrg0DxTUbJ
VEUhwQIr88vghSIyCItcPUn0JLt+7tkiQyvRQpUVNfToj8Y0x+5IhSc4G+ZHbEyg
YNstQtxrcj9D3nvpg21yW2/mHy5EXOYiLTW5Z9h9aIO4pz3luK3G4uuqQj22DYpV
zOXKXb2S6dzGP5FDpvD2fN++1DUGTg7q6uUbcAcvbVxlv/KNwdE/ozLjyqC4XHBm
GgpQAo5IEa9de1SukO5RQ4m4/3tYQalpUg9s/DIwPXzgnF/0WQeb7QyruoIQJ2gd
nw/+0yMmmdsvlTEJKNvvjNRVpHTsdrAT2FQbOJUe6bOV509qPbYpKUsBWZmfSUhY
sm5n1JJHh84LPhtOCqd/RG0bC3MHOLYFgg2rUluguy+q+sMMjvuH/ZTzTitAYSFJ
adLT65/eSIAKskrQwNFpDppy6N4gHTON7/HeltRCtvR6xbq3UODYBh2Ae5j+syuA
mdks0BEPWAcTg7LrfHRUSD2dHlpKr20HLI3h9Z8P+UrFUy4E9Xr9J+AOGmRvCMaJ
mzLHNrkooMIVr3GvK78KJ1oh9TCd1kZADS+/b145WIxMpLAhorMjOBDUzmjf3UOA
EmzQI66gPSK1Tmwb19ZfBC9ROBkEEIBHvKLp1tyJzUYoOcoOtEfPa4dmqqaEGVfa
bql5Cnqz7WYKpCUI4tZMwXJ6cvqNGBx2ahEGwdSV4PXg0in+Zz0ZREZInP+IHISv
NNeR37v0CAyXKmhmf953YGgX9jjoC8/CUdiIeCY6mfqJcGcJ9ykVrH1qBJqzIcdR
IoPAs4DU28oQe/cs9yhflOfVjxNzVS8q9+FzWbinBo38r2kLCKQ9KwNGNyme5KlO
0IwK8rn/C3/JJSDZOkzvrEM1IaOM1DD/1DLJEu/GGKW8gs2Q20dCwwYBvk7QCM2U
shKF/fyHwX/aDLuXnaFiEBQlYJIYfeY8zE1sJ9N4TQ6VN0L/vpV3lDk+VVd+bkHe
ZiVW++tGd5uciAL+CD0NyJuqqfNQRyDCJTERphsPR34AtlUQy/Tf26c+EVNPeft5
MNiB4sEUtHs+tRC81Ux9ylPBCduEQbeHzdKjwOKdgsMETMzZfDCOCD0YYF6hiSSy
K8TRMEuF4kcddm4x7sHFQUqRWqwf9PPIwkbKdIDVitbWHX91Iut5N+aNP8yAXrVX
MIx7CE4yYO5oeKou7DAJGU1s9Ni60cVOV4CYAB1zWGKSJlKeKgO4F0pYZDCvL0Nb
i6SvRVpf5SwKjjNdcO/QPE/6y5X4h9xW9PjpyRe5LZQW00hRe7kw6C7ij1DbobM3
gPj95P2ZPkxHKns9clOy9P5ZUs0fX2tPK3CBan+AgxS8wOlpLB9KRbBOYy13exQJ
tIAfT28plL+fd6Pc6ZY+VkFT4aKPMeFqsvdykwDEG195F85a3nVpBGeC5zNxFIzg
Qmut4NKyT8rxH15fxxIw+JFDu4rEt24cJOLLkTUGPpUPoEjmtPFq0S9JeKJuSUmV
RREvftoLFcQEklHh3sxW3Sahpz05vCnlj9djEXQzlwgya59TfrYfCOuYy2qlkNom
RnOeawl3Ux7MLZw8LX+TTx7fepKp52DPaAFmZ+5Zsr2XO1t/lV+bk8WEiK+Tg4Ez
7XPApidAQeK4Ms14Gykfc/Peo6La13DDvIZCHRYcCGtxqDYtj+u3EJhrwe0/NRp8
ivhikTFXVMqpwdbo1cpXReWuxm7eSLEhgstfUJU09acGgEceUxaM3pselYiN4V6S
jkdJLi+nxTgRIwYSveSCN1H7RaLm/vEawSI3dUDEnoUHBDAsqPjP9ep936ghTrG3
PcwjwIXQnHN+qOgvNyzaQsgg87Bk862btp27NqSc5Ibk5NoPndEMyBX7PrG/Yhqe
Cqb+Pi4zpaVKLe1u+zsmLI73c3fAPYnbk3313917I102faxGiw5Yg8UKAmzVzKd0
Zg6mPgir2Kj6HLoRQMG5n4S9u+7VwCYJBvN/U7Iva/m2y5bA4d+xp3xu+Fu/yQue
zbfCnKqDrjv4b+LsjUYKSaK3Bnit5kzinMbR4IGGrFKPdtm37jV8NghizuN8IT1I
T4YuJ2BPOv6o7hExNYmH55Ny6LNk5C8I2dqms0pAVETkV9rQHVLyVBbtT6on0wZ4
uoA/McQuExOSkWEVxfrR1RJJDd0UpnVe7UDpiFVP9YkjJrdYHUY3darMguKo8pxF
jo4O+gGOTEd4ssPuLmvfYUSEDWGZJs8fyo81qkDPP2ZQ9G4/8x1tm+ZSpsxdPY5A
24ZTfXWbmeWOI/+vXcMYfBNJaYilSj74dHGlEUwWM24dkzNd58XDCpFW7xinfqom
0B5AUuQK9peR+S/9ShKFC16/YoJ8ctz/zYXYbfjTw4ZUvd8gAlzCh0MbLtoSHwxS
l15iW2Ehg9t74qzpjrVLiKxerbYWZlclePkw4cj0W3VjQW+kVAsq8ElEOPY1cRsj
/FifTw+cfbTpE8gK/Dk1PEcp4pYshQbftNRieQXmPePDZtXwoYY6e+MlS73q8831
dRsX6Ung3LGYHw9FTiBs74FqhmE6/stc+emNwDdz7UWEnVlkg21/tt4az87wS8+B
+yU0o4rQWVWLhZKP0bVhncjQ16JwRz0Y3dKZiCGOw2dbRd/vPoIV33JQahl2BPuT
vdxlZQ5CW5MwxSzAWXbkVVVfWbO7gekzL01trUkuVOg0/NL1kkMVrAHgqEt7fAKT
0pH8gwCr8lNIpOCfR8jxaAKyfZLESQT2P64zdki5EahTCOrrFxT3nWa2on1iiUD7
SY+qCp9llZ+vWjICe9ZsBPiFgMRtEHRWlc47Jjdu4L65WciKneBZvtcPGTX/q+rW
+PgWMm60OEstsUzU03QwTREFrGLaBwqGnqzj/G6d/KtBK6KJD0ubbiVPDASV9p/s
c/r/yjK/vYsdOMcYOQE6SiSpHw0zT6zkfa253zYGUofR+nYsgy7N7bSt2KevP5CS
RpcC6MutgmsfR2ueJhJbEfvqi0EZyhUFdEfSAkuCIzTWKV9/4okqZc4k6AwyVJ+w
fKMeT0eGAJbR6LiUK/CGSlxgrwPCVSsS83nR7AMtaxnSmtsJkcRtw+rwhSVYazW+
pLpCuaoWhZWeYng/k/0VjpCRp/9O1LuiRzvvUJ/Z8DpgVLbTU0IRs2Fgp5pOTnye
PgvyelFk05ZA7V+tRNBiPP5DGnY469WW4z76sS58YZemVoeE2dBPbOXhrpUi66az
jGGtlSrDQ0MOpOYk2cjtXN4y4mpPo2YEG0l3JLctsm/kEf1hFF4AaA4c4G6eClXI
veH6dhTjQGji3Q4FK2JjNczZVCdEudHq+AeFqr9kdiQGtsfYA9EnIxoR7XywDM7n
QjqU+QYrQdnpaRQ2uO/nDOo7A5U4VHGFrycnnTyGttCx/7UkYGIKmxTunq9f857s
3/i5v9R0TYquhLjHtxOdUg7+NzJz7NAJgaohP0fFbr6B4hWB3j327R7a0UQse3Jn
ay2fB3EHJLt33eErheDHNX3gxcwy/f+3wXrCjWqoJeb9Zuyck8l7La2ClMhHEPOG
RfFXlt3Mve0sy4ky63JAZSZyqqEj97BNPKAH8EftFYEvv5ON7DtCFbg6Fxe1D2BS
QiRY3aSmkOSXHM09vZbO32hpnAq0w5VC/PfzHljbUUe7K6Si/UozcGHt7XZN30gC
VLHHR8kHnHj45arELX9TBu74Ou70Us22HlfdhtkNZvfDbFIz/0QEipqsbFPgWsNl
+ESNjOhL83pXMWDUvf7N2P7Bo4ODkz4J0rkBbxqdUjBLmNkHCXot6M61c/hsS2kG
G81LavbBzl+j4YaJHxMklLxcAziqbzsT3qUoBsO2RAKiEH+4UQdDLobgsXJEMYjP
4BLTDrCmYNwLCYRkAHz+ISzGxcD8RhMax65STADjc8q7/VvBIhtbg/bypq/URRhM
GJ26ajatTrzMKHp5X8SLhNPlclxqGy19sAXdK5MNOkuzbhg5CjgnhOPlMcJuO5PZ
fUEHJX4CIDpBHEbIoIS3YryVm/VHyzu7fj41n1r8qVDALH3ek0LDjNamOsef4pIH
eWqgv8cTw0ZefRvzwr61iu8kX6VZoBAFKQ0m+ysqZ/1i2NW8IutZcNCUqTJbkGPp
RT8iIFB47zPZvoztui17DcWbfYkzCrwwGotO/H3vMJavz1IPGhC31wC/UtXvx06S
oaPq3FBVTa7+mJ5tPrkbg6/VYNSwYNnbf2uaQLAyFQ2x7X6y8CPKl9gUuSLYZquy
2EjWgmiKY404i2HECKLKyksZ52+9hV17IS7XFFzsD2vVnfbd98TBGat1AzTYDwRa
tkcUcWF/3OOC3yDccTPO2jNv6u4hbvOfjumqiq6Z3mwqVSKPlstuQUfAXxXplyGy
qjNFqimWT1bsgHQV+WUr1k5lNL0EZV7Swb6eajworzPmLExOL3KEktskVNUr+B/g
lxAfDkRFBCGiS9cNxbBd1erK2Bn2zyfehIQywYzcsoNook3oKUgmlxSKiLy4OnhR
LMM5FJw8ztuJhDkqx8yJtQQzALNV0RSy8512ox8Ok881X35jDnPthaEUQcqwwAwN
tS+twTz6q18ycUU7VUBhaYbd9koqcxyn2zZ79wb89KRCTYO7ge3UsuYDTIYMgZxg
hossJuGntoEyY1ocKFmTx9tQSYZS7dGLHw6r68+6COcfBkY8v1B3F/9TNpAEo+d1
cVw/GJKsS8kvQTknpF8mf+SnOOOuZTRCdHseC35eIp41L50lqbLakvLE7NRGoawp
Q23sYuYah9O4MBMelqHWRi49J8oUQsIwSqut5DD/WIiHPTcswWVV0nL5qLeRQiYJ
rUda4UcLKLuSO2lQm6zqdXIkYwIQxMWCrZ9cdRYk7V+ULmyx3uAO9dhZLP+hup93
W35U8+Lbn3EUDh/HZMvTSn/F3+mEAV10fqpXAAMb6Tgh494FyvrA9jCy2risuHdr
5ZV7csgN2q4gQP14/G3vPy4I4VEIoiK1sN4hf4c02ltm1cjHHSDP/vkMR/Xx0GQz
oGOEHnK6r+oIk9HIhbmWWDk5xlw0B8nAUO9qk+/8fZijhFR9/o7UgRszEfy29jCS
eBqLytaq4jgqbpvJ/1PT+Ugldyc9L2ZGd+8a4CZ7/X+Bq+XXi5jHNadL3fiInlH3
pBAfhrxHoFaG+jbiE1gn6EDH4UVGP6i5UBlxR4Uho209ogjKWy0Vxd4qOo253FOD
trV4lpmvEkLM1217TBhzQKXAzfu6TReM70TXyaZtUPsaN1APvL/MfvJEJVBvTTEC
YnWJ6V1x7Yfy2tU2oHgkP+k7RW9/Q3CgZks798cDohmORjcxQGdthxIs4WRP+gJ2
Dl9MbMAmyt/SteCViRQhWCuNZ0dGWHJ72WK2s68USN0aic9UE0aoaa6QqJuGNO/M
sp4m+ZuWCJGAJHfOFiSz9HfVXhHnFR/ZIFX5TMgUtN29+KXSrCKBo3VdWA9wvsKP
oUOgkUbMjl6rDgaI6zpdIEMUlMFuDyPE5/s/5SWVsU46WOSy8tF1peFdQ0eXdGpO
5rmEjBwJ4ofyotcDXa+XFkD0cqi4FPtFO+NZBVF5vy2CLmtvGxpKuiDn6+p0e1pQ
h+xQpsDZj5i5DWGUm99vexN5wITn92omk1/jreTIQNsErRz4T0ruPoK7vcXdS/ic
YLQZ4NCMU/Vry0aLtUtcWu8hI7ZGFILm84EUF/8Sg7s=
`pragma protect end_protected

`endif // `ifndef _VSL_MSB_SV_


