//----------------------------------------------------------------------
/**
 * @file vf_reg.sv
 * @brief Defines VF register base class.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_REG_SV_
`define _VF_REG_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
feUgvnfrN8nRyaqhuqQqAesRI0Kj+OFArm6mI9o05Z0/M2nmdKe6qM+968tuyb8z
1852bjc0S0tTG1T0hSq4WtHMILznxEX+vHQMe2VMa+nYQJqnCzZH1BfW+vjFvGDi
OQ7jjlgx4IAUOrMFmkA0CUlwMthk7yVIPuoTDUUtXxnmq31dGIYGDpZAOj5BHHDM
nqrqQFDf+LrLQZ5qK5d8qNLAA/18URm8hIyQ6VNi7j53sBEHvieNI3uWsyuhlCvL
XjnAdw3xEuQhpJv4RBIi3D10sAurpPLJFWO3Jqbtq7k2J+t5YPYZv0CvQTbkIhLU
o0VXPEopdx/f10JYW7m9ow==
`pragma protect data_block
ZLmvqZQbulUT37Bjve5E+gYmJfSl6JsQrRh5TJhanBS2mIt08aZET0XvHZm4cGPI
9nPQTZ9Q5rtVvP3ja07bJ6ADSMymGzjfywxF8ocJYWPYy0NutHGgajmj2j27hNww
nJXh5IsNqp5dmnGY07SlveTP3S/d02UDP/XHYccsnb7tVn0DGsVN3LWdIsNEW8aE
c0unP7xnq5Vz3bpmM0jkTtSfLNNlAtO66axmku+AMyrhdOFVmuBz1vDKtAi+7FU9
OZOACMtVGaNVIroNGBpcVNwkC+n/qHX+/AkDF8JaCVlWgpY5OCyqt+ry6tNGKyV9
qWyj40ncxKG8g4WvwKASxpCPPZdtJKbrrKio1hvBAQrQnh7k9DZ/n8bBv4XwGAEq
TOyqrfksuE6zGh7M6FbVJGO9ExepKrUMVhYyXfEo76k6F9NDezZNl7SSJBg9v81Z
wyc+Y4UG+N2SEZsAF2BXrO9FSlPAYswJu/TMij9v1mqntfM9gkFCqod4WTlNv232
0MYeZRgfM20yy0KjcMAG72vzvomJPXIMaa214iE/0aLpk+7L13ZSzppqte5K90WE
G9aE+y4aoVadsA1AJiIiWjr5KewlyUTSNNyUfxWs84qaDTO8DDO8GdySvYOZARvs
4awTVX8lhg1sUp80tm/2jq/zB33cBMW99V9XcKvRldEXQ9/Z84pMz4CnLUzpPLgV
3SPcgZblVxeY83IxG9Hy5EU3OdP0amqlKIx8zI6dlH1xpjyyfqtuM45qJ3ZClu/T
epfGhsNzML6CFxuO48oxi3QUKuvIsYuS0BXMJlR/MulD6QfkqK50je9cA79HUIa7
3OuHS0B+TBZjqO3haa4wBDdjLzVJhmlLDv+prOoKnD4PsI+q8yKQ59csGkskotmz
J25mMuw0GctUOrrDbM3iRyt7XV2jv9SAiBoe5I0TzgOqFSqVXOx1z9pyxUhRziYF
XRfgC8Np3IYp9RGxeBcShFocSwRIKVVsbcmGl7T8y9N481dilZjrTUYkg6GBsDJo
gc0HfGjfEYhjF5YVo1tXPTmDOxLL1BlEg0J03Hk1CzFuhCgiuEvct5R2/grIlpP7
pFfNmvBHdA3Z7udBziDtTj+hkb4155cvgGTLG3XtyVuRcQ8v99t6g2ZIlavCYvLb
B/Hvs4uH0iejw7tjOVmp5LuvPmEovHCj35tXKhkh8Y8aK0640pWOhC2yhn7Qy+1d
LCn9Bx4TA1dxJqf5cwSU7ywpe8LeaCwIh/4i8ZG5D2kyBpj1bHdyP0Ihlxlyb51l
qilrl3yFd+RYMI7ftSsiU9/nB8Jg5jKvyK9C+3PbRn+4qeb2kMg1YQihZJw5THak
DQ/8dm+hJh1ib7gB/BgYLBnzyyAA1tVKh6n4cw3p/Ob1MWf10hps1DQG3bFALBck
5iNCFcpJnluRoVLkBp0VL5xoBpTzuUgbgJzuyejVHpbFffnRcGHs7EQIKOUSJrGq
HJxkESanJKryu1fEw6NvVHkDhIAFILWlZqKcm3BaMgUQrF7i4NR0Tn752/H72Ysn
/YJR9wYPWoTED4WB841DVDFUI13ORBFryndOhqITArPH+XFu1R7UKADV3ovwN+gp
UAzLe9qwdHT448dvhmkBnodpm8y35K82ZOAY8QJE3QSY6R93iEBZDwhkizZV0i6Y
/LHsCCbIcgpu79JKtvltKgWMqG6oOJt3/w0bDqKrVkIzWid+zUCTDO06rs+4Czem
7n+mSQUtryfx8i2CNxkCCk9DrJOql1PNrunr8ct7QPhp8DfODz9zDE5RdqW5LLGv
0xs/qgzZ37F5rsy+GewrJX1WdwYDFDDvixd+iDgPuw2LVbCQtERvlH9c5fRE6D6S
dcREgPlmEoSDXpm/KrCC9ufSJprgPBj7B5Wxdpzk/Se/g/GWgY4fw6oABq807T1G
N5Ix5dtBYBg0KHFRUgwGr8vl/tg/wX8kaSutOr0N6mdKjGKh+/os8iM3BQsUlEB2
b3QkPdMnGZ05sSkpCcQjbO2+cKJhG/EwiYwJk5a81vRAWNk9Yqkz6hc+JJPfHAZp
iym1p4xWytMzuRqxQxXGNTcwb51r62nZw6XUUkW2wALFs3AKQrUMbzSXEsfMRGjC
F8EORXKkEtD2usoaG0p3uXhJft5oKcGwvU1GxCjV1qiaBQzEgMfVHkpF0HDh8Gkm
g7VKiMIr6EYRhq7JKHbKg48C5Qoxn+nHe87/EURdmpguz1OXva5K5FJdLR+B/Hpi
vjsZE9u7kNFEFpRuYr+kxvvs4oFEPAwh54rGAKBuujxJ2uWng1spaMCKd2HB7/6K
9v6VCxJIBBBU7EBqi4WmI6+Z9Y1VzgHn2dJXxt+S1mPBcOHCqSP+QZjtHJ27eBuw
nkF/e2C6fw9VbGLvjIc4KEHg6PXy8rqVJ41BmYN//ZL1seTLjilQV/YuDkgr7bng
P052FmDV50TZsYvhQjpZTJZsGQzkVJwtA0PFXL12RcyZLg00WgwSciXoWLj0iXKh
45r5oKcMohDvT07YPguM1c463eBhGRNvedvL+lo13LwUBEmNRl/DPOdLjIsR8NHK
JlsdnW9aUJB9ul3xEREt8ZRbnKL88esjeq2WEsCTmCKiy32c4DOGNoRNUCH7u/iq
rfsjjT4I09uayJJDoiJIp4lzPBS/rGFg2oDztnwRPA/KFbXCw/8GowmNwzmBKctS
4jBEDw9jS9Vxqskz4AmyCpR4IEmZtg5pGPBNpT1nON98pcZgcPdYzPZIbbfVwqxf
c80lzY4AR54fWIK7wizjhoAQDSUKA4s7zIdBRQW64F8QjhYHGVQPng7Aza/XCFBc
q0rfOYTumtoeAgX5kA/luIeDSUApsgtw34g0SGvK0pfG3cQK8mVfIuHOfSGgPPwp
XljN7z3FO5DE8PStmNmt4VVN12OULioz8QBaUqwQSUq5qOY16V1CC/jrKS1gPh3D
/0N38gq0j9dRJVICoNc8p7oT94KSliHaNhJeDU7GhDid5oElUxsG3TO6QU03dUby
vJfuusAcs1FMmGQ3bQvJYF87ibph01GZsHFdwn6rEMTyqqBCibW57wlarg1ZhESd
Hi0d9lrTbxXZus0a5sD+/sikAVE+n68EoLplkQcjNDh2GHMvgstd7ZfNXMjscpl+
oaDlbybv1br39x5IbQwsZrr0phb8ZKjkVr98HDLLUHQeo2l9fxIzqXbqWPzNzZqz
/FjOCPh34KsyDzv7fiYFeGePg9i9P7NmMd24nn433MNQ38ZzeVvvtJtSC/ptlxDj
Z/QfyTWieZOsIY5lK232mFs74escDHCtG+Ewvo/M6pmXeZwfZShQhM5UwGeNkADg
e0Du+3DFCVxbvvJMgo34dPY/rqb95qUNq1Amrp0A7Zs3irFfxX2175TDxhUkQJCE
O6CD12H3Os7Cgvb2zjuBKBresXHOCkvfrGIHBPAEN4/js/OiqtNtYcVpuo2qUjnk
37V4PnK8aF5JeV1N0Hpn6wfP6sVWwyvArMVnpMgN+ZjnBvytRhfrhETuGHsA30Em
Ji778QN6S4p3CuRrY8YOSQA9viV+DW6ho/nfxqcM3Ngu3N8MKRJJFJfRlaaXC2/p
pJpGWt666S59VEYik1skubKmhAgjWZGmA5se6NNk2vm1Je5Ur+3/T4Avr1ibo6sL
7ANGNtxXh21U0oohQuE3NPKzIkgHJ5gnQ/NzFJobHaxTUhHiaZEIAc1CgvABq+Pm
3wfUt7XH5lVQ8QehvwNRFTqh0s2m/auxYtA9GPTseeWAn6l+idHl0OEdyC97FzGq
UgLf3sBGwhXxutpA0TL+3IlXw13gwvKn+bnV9F2wv0P2xLIgR2oU/9vk7PLNDMQo
IipTUBN0DAIDc0CbuSL3vrbw/BfO4zrwuv+s+dMTnw5dPnKlWZCspPMb47fukY25
IRBHQ5oEzuRIq2k7GQyHbztirOKbnUvhEXfe19QgtIZlhtcsSiwmFaF2kuvArWxy
+JKMvuH4HWXk5nOXWz5LWT31IGZdKk/sCp39nrjWomeIVVB9RGzoBcNktA70ZTJ8
xYv3hp76z/FuuZUzfb+SJoJWk2t8Vt5LMmKfDS3jf/xeCrA+0Tbu2zHjvMo3b21V
x9FDYXyQRyQR2+0nPTi7Oa7rdVB1HE7bdKp7RK5cHOthbVFoYMBQ5Z9xqcZSo39I
7VJB3UaenRfgk3SsDJufaon0V+yBH34uF9yiv/o7NaRQgBHIRNI9gbCY//qdTUZK
j86GHJJdomp4GtzpvnrE+XUuEHvpIzpM0RKsFuhZA/pDApwUHh4HzKtgZzRtMlPr
XAbE1CawOkhqdZaKK9R5md2UXL0Ard5vH/CamN4Twpyom075yhpIxn+XY6hJrClG
QQQ8mMpFQbAq4cJickYD2BvlmFh8tQE/dvvP9QBhDSag85XTnqQx6kdoL/v2q+AI
5pQRY5XxSm9S+3wvHihqQDXXZiS3VlLLQxhomNEOT5us5tWgVFw1KojZi0ddzSko
NS8VkTNN0/1/YOenXteC9vKqKXngXq0O7ovAGxedNaC167qumPBpPlJP+RjzcxUA
119M7R/VD2v9By66YP6LjqXLFZnGT5hBSwdWQ7HaPfdySkhoShfwzvWLpWTnxsKZ
Tf6Kndt8lNxrxylHDzAriKFsLTAz6VPy9Qkni5d2dS/KzChoPO7gnNen2n08mp3G
Vnoepv+fh8y7xUQ9+kUuldhbyVoJfBxJl2Qs/6bbm/AnfVxOPgmY7gYXnQpUyh1v
T6ya7j0ABve0WGIxypCpYvhPaXexPA3E/rxlmmT0WouMfOxNXfMZMxpHUd1mV3ua
ShnGma7Yt3YPhzSY7Hvn7/Ry7nltJ1Mp1pNESGFvDkgQFN2bgXQrl/2WQWcVvisc
DQ/kk2VWq8YjDQJHDdARmmFm+yPeKecRecTZoJrwLAjMxQr+Q14twEEszHK5A6uy
x8IUdEtsOXJ44CLjr+NRsrO4bvHwqTNyZCHf8jtUdcshEaipGC8tW8fLmiGL82MJ
W7TCX/uEwH3spWhfvBnpWUJ48aHD5990C7/pJSvVMZiK43rjDQf2/x4k3DGGRDqi
YQWhL8B2sCaEcuLU4CuX4xgfnAImmHnAdqPuTQB+aSNbKTR+lWCAuKHZtTjBpQdQ
OgVSOq5bI20TmycnOsLzB2gGAgjSLBAoNl1byllMkmRbBhCZTuEKA+H5VqDqv/lr
oY2GLDOwyb65t4qx1riZ2ii63hq6EcIK+hlRuL+Yu359RgTA4at6x3FJeGvHeLcG
AjSpgwnq7DpzqNCtgylTW48MLyYhZQx0fx/aEJ8s/IroSWjOiFI2KIxXYUPgJoGw
9URHK2qJbHS1KA5MSipLcKbOcaOrMgrVghH2M3l4uUwhI+PD+ixUMVyRM98CRf82
Kid6aYGGnHam71PvAMLNr7WzRQRLHq6m0KEdi5PNT3miMjR4ZknpxZPmYvWGMdnz
0bWEGDo80qSGTCHMimRHtu1gRCnmzoSMqjK3ivxeiY2exeoYoG+rF1/BfsvQekC+
B2bJ+rSAZereADbf+xDRoY6Ig8gT0Xpac9B+Ip9TFZxdepaHBkKISi6gve4XNb79
jjivQb5Ba+M80hIeQbqwSzWLHi+IBB6wpAJzjh6x7wbk7zPBzv6jARYuSpd4YxTe
/eQ7ascLNFcxyu0oGurmnKD8IYUz0wJQQV0yjcPJhtM2rCmoAqJlE7+/tz9G+4EW
GT79wpnhDYnVCD0h1LCAmuTPYeygTuMepj6Y8TIgxbQe5JPKkuTitMFQJAfLjqlF
0kJM2XU7Xp95y4/E2kCm2KtrPkR+gwh+ORFv+1Wk3ogtqguvrS657D2W4q2iuYmD
54gcrUVeTx464738sPWtkx22hIUMSWmMldWglSKKR8XHxt9dDwGIf+1RKPhQWIQE
HLxNa9KZycuahsfS3oVj4m7jqSZ/Q/Avs2PbTQGM5I99YCs3pyx7kB6RDIDlLCqI
c8hJjs59pvbHdba3ouJ0HrqD5v/2wRlayWocCYpOXRZ1++d+F0nVTjzkOkNjbvZs
aiqq4PcBiTpmz7r3NybSkmELrBJqPwDS1iFjfqv43yhS9erPWAsTdiYEtuGI/cAt
Lbo23MVtCT9gog9tTU8iCymE+ueUESI9str2qTsZTi17CWcNEQg7FCjEnB11blMQ
H75OrP0MYfb8Fkd/65rTdhUL/MOZi23fpTYO+cq+brU7i4BSWErXqxAU0lhyGOpF
elaVG8NPbdnb0RpKIgxncLevpHXhTsIAcCHu8FWleV6FXC5QltfBeVK4QPSPRHCB
pbO9pJnpcsBBzowgmPfNuFgWUoU+v5r7Nij2SMMfodabOUaDZoVlHCeLYX+hbxti
843ECOrUcHovrg2b/jAqKRFIBX3T+WGOeDmPa8WnOml77QriQopelein26HOjQfw
2C8jFk+1IIpqWtKZ2Q9dri3e+ZrZIrmz8Gpe1fx/gdcaDMuHOwobTu6M4IeC3uFz
bDLT8dcrNU+c1hysGgHE521F7piwx8ICVy1nGIOMg7hXz6FS1lJ7A6Y7WJ81SSLR
KC4JeAzdchoe+yQ1HOBf0bK1fIYNTzQjImbTsiU9HA9lCalkcf3VKOwVrXPICgVc
ekRU8j5MUVujAEl291RJkQVfzu8FV59sc2sI8LYamQNuyDSmQ6kYNGhE16/cxVNx
5H/wi+QZ/7njdE+li54/tQgl/k8LosvCHjokeDvkp1Y3YVfn5H0rQS5KmAtTyfaB
2JgkIC/bxsQ7CcBBVW40diNzt39GT/+sVaqUF93OKjhrXNT9XhC/w/B7tY0fK/5p
UaQW328LGCK6VMZ20d2v9H1SIF49Vwr3ZnrE49ocCT4oDeAnJBQTsAfwnjODDKnp
LksTzA6OJ32bFL/asnR+yZqDF9sfkw3WFcaa7vC/w+q+ZcEwwcrnSAbIWz0PCaMF
Jh0WGgQt8q6fAllAWLrO0kjjRW6Kr3Yh0F1wc4JfHgMwH/iTS4N9/C+6MXloDx2y
9AWwWoPJSNNq+4lmOeAWmoINfHWoRuiUfrE76o+hJSaVWOSxD6ZzI8MSHF8EC1XM
QL1l0ZXSqYGwCzXVBBntRNey+gAxYZY2InUf/IfB+HwL7uAeBJnqZCJ8kk39PhJm
OAPxtPvtTthyS6l4SMyL/w3uXvlErqEAVU76rgT+Rh80R0wrsIAdoSGgp1rNWDpl
OOHQiwQJAZ+tXVCR3VE+pXUz+I5dI67C5RmHuYfqiYmac8dGi9QyfKk5WxAhyQF5
38ZakFkRwb7o1kEgR2CdMKq1psCYQdB/0gHAtWnLlxlwlW3BpO6gWt/U1WTXFJfp
9gx2O+JEh4qaM1wfNF/dsTuqx2V4B7Prj60msTDK7LVxjbpo7y90UxfrZHZeg6++
54V0UxnLA6gLH/nO6WO53iEv3sCYe2B0bh362gYkoqz710zpCpHAbBHVq0rnICXV
//4tsaqYzjgUfnIO2kdL/JgvIKnQkeL/MwoVk6LkBIwXZr1OVNwRW8Gw2LACcrVp
p9j3a1nfbTyy9d5YSaKSPLd4BZGi0WEMkvewkgVjdMz9FIWupnkQKc+7nuEznx25
J9nCeZlaroK9b9hmm5ZRMnw0roDpsVt6fJ/+XPjwjYTIHQJSTFgQp2ge/Vv2oFQr
uN3WzR0BXR9fRkhhiI59E5HAGoPIzU32OSrQGyuKF6meYL7nk9vKhY662GJPNq21
U3rCm5aY3vvqpqZJUGZ0ygjUwOwsFt1djWZNnHs9pQy8crn3cKe9y7DT1fXm9XcV
Z5auQ+iN3+pyqIps6l4zfak8F1LqoX/j2h9W8GOb3lEetRywvWQBkc+V2ISPdvTk
t3RS285quZ9Q2wFKmz29c3YId9Yl2Yu/bEJeiJDxWTTHmgfFEKefK4lC3ChCpAEA
VrPPscIdJ4r01KP0Oji7zHW58kIn/c1HkPjDv0mAHaj1E0GzOhx9unrd5T2kO7Jj
M8ejjJTWEY2UVxxddWoRnlcjw9t7MwitCnfepGWFOmJnOFKmEsA5xhcH7UnMgIwh
TGPUi1+Y+uevaYK+kX7s/pOpPytxg83dEUmKJp1ojGFHWNJHRzwTgZBNdDi93Ipe
UV7UbTi6iQEIqOoLbRSSXTY/14QdwqatwZgJzm4u/6h3mU+uLpRgIX2+QtwtO5qS
V74ZbDySpZKeAyXIEjypwbqq9Kz9B/A/y9rk0Ssg6m1YcnUgg2WYMbxeHvy18rYd
Pj4D2GfOn1q20oIwH5xgPrTSNFutyxcQ0WvhhQeKqQVMrDZHGmGiUp0fe+1F+UWy
ScFTkrDiWvUe9x78UhGuJTcz71xSsuJn/d894ea0LJbQYLWIZPddAYVYYpO9q2OK
8wXIrRDeTpdkZQ+CoBRb+Um4eEh1o35BxFhzBuYAwf1Pr43Jqi48BAXxYqN/mNYw
uMBNUE7YoEJQMffIz9IhoWpni3vYqOBAj7/ZXKztIGyug4qWLRx1RS0NTy2JtYWa
VwEjBniiKT4loMSgLedsTenJOrJuiruNrtcDyLrozlT5KHkaeQfMgqoMvxzhliGm
/6p0vLwKs63YRpLgzMfyW9JG3oscgIsRdaK4pZDZ1LUdBTRA6iWj+nWjH50WzOI2
FtyJWN/6Pfy56TT+q++ZNrayr7UbZaoRTyEFXEiBQkMWs9je9NZ9Vcvuf5/X5ew8
RHKTdmxoQSo8IVjpS28Xx2sLgC1YniDCPuTM2q+tQaFAGXeO1Y8edIgs1B3tgGqH
n2/aHQxFlB0OnqwMB6SCggvYSMAItTzx8EM4quiN+I1ShptxI6vYpud+0enVK6Cw
XYLr99WnWRv8gGbIvJ1G2RnleE18byrjeusgzeiCGFyL5JjdPlMAzfwfc9y8MEp8
ng5P4Mw1WThGdECFYF+NC3c/pkcq2SpyxIFh4aGYdluU8iEakOrhrKML6LMSxDxF
VbMOKnGmuGmBK2nrwGeoIHv5lZIYvt7nwg6045QuyMo4xWpiRgN8xk72NYgFBy/V
Km0IznPIFQqDOf/dJr3cpNY5o9tyxkxd54XUndhnVV+sXUQ4rlpaIMpr3aBFCplo
zq15oFrwp1SSxqwUcpdmkBJimoeEvBO3rTJ9pf3tLbGY933TtT6MG1ONrX/KJvBh
1/D6wn6wLYt35nuWhZP80DHidhbSPJJduAUxEBBYTYRZj4SPlUn7UhPpwUFBqDPF
eb5rjazJdifyBMmBLJOThvEJSoqFOxGGpWvh4VHSS1zOA0KrYwalR8feBmWvSqlB
Z1G/mayg7OGQmy2Re/ZQFpL+BMOlotRmYq+zunERfnsV1IzOlDahl2EvLRtQNzX6
p/668lFbGMhgR3mrgiJUuImqpS4E9Uz8mIzbUe6EPjlng2if14sVCl2MbTm++yXH
FX0MET+l0YtbSYTXWXaSEmOwAsptVEgEU6z4sVGE8XTrhz1aPNHRxxmL1xYmI+5c
OG71EvBAgWcDs5nKCUunXudM561VWXw1j2YoWCOlJv2Q3pvmYYGZLmjqVcov6Xuc
ZA3e1CTunez+2NaXZUJqUcxDgaOSz7ac2/i0bD+4Tl0mjXlyeMCIvVyuE2K9C/pW
B/mmBAKCllyPfHeBSvhBCsZiP4cWsJ62zaS5u5fOEFTz8ECc7ZGwA+hnNKVwYZOe
RrDpcuPCS2RP4hR1fDwiE4pDNpa8/K1gacBTYkjF1jxCwFbDayzLwo//5+jaKE/4
JR70lPdM8ynDzSumytHKgY2t5BO4Ebx9Y3ga5ozIX11D0pEn//CWUx5XBryshqWZ
sSmRQnnzUQk8jq4jJh1v2OUbuiyqAirE5VdbrVBeUSFC0k4sJrH5rvbpkv//tib3
YQbrVIJjEUWdXhySeV7kLX2m9ZckTnP8glkTQzWq6/YcxpbygJYdcR65PyxEJ2yo
nLCrofShWNh7wj6sI2iOl7GqfnPV6AMimCH+CssR2DjVL63tF900y0GhLNT6ToBm
PO/zZd/Q/bytFkZ99gUVVPKMjRpdWB46TLWS4MPxC29V8FZKRMvTl+QsTKOpMKWZ
BJOr2Q5kXuptRPmKhG9HK1hqyk5rbJs33JCbmUNA7PXcq9YTgOFex9QJu1f/hYmn
MeCMkf5UZc5a7ryfA+/HwlSRSUeci3dCjMViZ2fvHfjfBdNkF9lBt4zrituJ/nVE
CurStfa9lKZepI4sqRNDVvEIDmvzPL+dP3UP9ryoGZjG4dsU+DSrfFRF7FGyWuo9
RDjpU648fX+54TF7AsaH2upgm9dYvozsAXwgek/t3vkF+vGcJ+3fVoSUxgZzDKpx
NxmCoMTbEXRuTvBS1DNTyDzxRkgYCE211L4iFaq+oUOI78Tj3W9tGxUbs5UWImR5
SyyCXEJrL8iFPM4jdJrHQi/ovSCQ+EGSk/mt5XhALAVedm++8b+5OYLEdeFAD8mr
yAU8xUMTSpc9+UNp9yx2xt+c3b3qQ465ZIFoYTneCz88xUah8BRu7sZGh2ajv9Vf
pmKhnjLBmFADMXcoSYvNO7tqLnJ5KBnnmXMg5BREqTK+gaXLa/XCf8DlVLFV7EGx
zmpm1pEQx+baBKIWzRHCC/UwYqIFQW6mIsIJJicsnWzIIVvAnPpUbb8siHchMmCV
r4awb+j7ZDobNXHXWuUzpOEiQlEQbN8OZZ097O8rqKC25dBgHPFwopeU1yf5CSS8
lgTaHmnmxDqoxJSadmTeLhFRLbwhVRbAN7QiwFQKcKPW/w0Ey/0kdp71oX8qLImW
WyHvZvf0jKP5XB/AXShAXL1knYF+r+jfkoUL3hlBAK0O37PAvKA2nC7ffhcD1+4I
NmVf9rgp2eTupzmxFwuM94+dceugso03llTnGgJ6ae78LnHkXSwhLMsj49Ht1HBd
h9KW3p3ihxGNPed4jgWPbOSGdECGc7EKePxU9GUv1cQR6lmN5ySB+64/xlvnlJ9T
V4NNCBfoxFoN7HXHlDXZUO50oNjjhygvmKJKlhmDBa8szlUOzrx16MHnU2E4MUSd
MXoLZFYebxLEOMfTjByXkpjK0/AD6lkr12mqw5YApK85qnN5T/N02LIWM2RkgPWu
uR9rzcaVZSbIK9kQPN/3rn+TeD9RIEJUYGaxVr/glHAB3A5CaQS/6O2KTUe7cCNU
Fz6MJJy/cRsc7oUFJHwXVaMFKeNY2qmAeKG0M73TPp3dSt44375IfDEH1n4eqVuN
TsOuzkkRrpqVZGe1tOC3+g/aH+yyWiAMqMTZotGoVLmme3THLzJiBZhQZkP7bZtC
v4f+g+vwRZ/iDgKTmwpzpjDIbb4ir96uB4Rwc3dOdj8dXAm0oPYbcQ0kG0XfY1Wr
bbhIhNkuOunzzvCMO2OLbP1FlTwHrxRTDQqdNxgYKTX6MZcMlR1EHRQCVaLIyQAQ
CS5LIVuI9RUlE5s/HDw/r62hJ6trKbdFAWv9z9+iEJH8/VViMcfXGQKl4+D3zl9v
wS0kOWnRJGdssSSVWIQLTXDsKTvQin6M+yg+a1H1jcc4GiSirXViMc6iVC40pLDV
2RXQCoKiMzEFLSSTeYhFXRf6XQxF25WwyMzfef3B27iggq6ppk817BW3Bxqrr3FC
khHxVwbm0HxWL5a5MOL6vp7zOJ8zv1f6+baxcb7ofCZIbKncugXIyC/vgKhWFw2I
YnDXtjboBAbbJ7x77RHli6vZMVnb6Vm6tTqwScJ0WBg6p1fKPf5kX6CyO8PfmHY8
2tpdKnPcCu2OZWbujLnj/1ve8p9mwr2TP+2IKIw3M/85QKPBfkdwqRxeqmSLfGTF
2j1F4Rj/Ypu7t2iC7yUDh6b78WQdHprcmugd4it00HFZ+9cBhoeOwGbnoDhNFL8s
0pH2E6lNQ3Pxf61FAeTuR+59DIm9gtD9mJqwI8k02pPg+mP0Z8WBrcMBrJaFGQlj
oN7SQLWtq1sE0CWqW0JR9HzifrgLsbM7zcxMlZcXzYCTYwTemfwjls2TVZoYTRJJ
IE2agfUGv/55NYrce4VupFTkHFC8HODgigiicsdOBi5+s3s8W88zumd0u4frevq/
wq/cBS+QekF/gTGTm7VwQj+wKe751O0R/BN0kCCVl9zDj0iDzKIz0+ieZVyhX/zn
OJAiy5n+wkkrvm9YvOAh2W6lr/alCLdgGe5ja+LINhfj6INuLH5qmsvXEycM1aAB
FnVXZ9MamicMgidFHvgOBFtAL/obbiMUAKQJPV/2no6QV3cpaQVH3Gv67fhSPojf
QeCn2yuCqYgGywsamIYXqfXiwXdX1x05hOgIE7fH2zXeD7l3ZEFf67NXMEiBWy82
ID8bnpephfy8Fi2427dcz922UoKlrp5pRXtS3eOxbZ/eUCpYzFQJM9knIAR/EkzM
EmuSGCIdGisCWBqgqBziJhbkim3Oim9Y1E7I5R6+57hDbmBWiBm64sI6QOQxJUa/
T2dKDNofykyZV2oUp+QFHUE/ZS2nFpDCtUK92wpBvXSGe05O8zl2kaMN7iT5aYqh
eAyVHw+QSggIS3woqB7wRboNWEZN/IOdmr5OSw+/Chga4KSesQSSZOK2APLlL9w+
7fLP7ozct393TtUgJmTBqZWK1f+zIuXLxGMinGQP/KLskNRjr8njxS4u9A2gQLTJ
IEu+3u8dv48zZYiGRr2b1jES+34JClVAC7hIW+jMTufL5P473/eGeaUUA8lNXeJf
x5Cqyqi+pkxEdLdGM1PB846x1bc0HhYGPbQCD0XUsqBlsvD9ONOR4LfJDfyVXmMq
ALBjIspJ6hYUFV1R9oYOrKmd/V8Wvc5NRIP9M4B/WzOis7/2TmaZm/GBCaDmTm5g
wfdYXCnkyUdzYwrCPG8oTqa4PgVGIooz55/BnoEDrtrPyQLaH6mBizDiC0yvW0ZR
XbYoKfX0JrOZYAVXsw43SRzFVEODnkEUMbESieIO7NZyIt6srOBPsTLc4a6lGvD+
1Li5DTZtkazJNQpoixXj45ryXBm4QQlDM9USqeCCiBTCKvilxh5guzzVNrYhngn/
EJSU7CBW/Zm6GqwNctZbeDs+JTvDBBxYwRMGAUJZ0n3qVGDCIdiXVUGHByM0esdB
mi5HhSGA5F2gU7aeMdfwy45ETcrVPt4GiMHEsgFNC1TyaXpo7EvGbC5Bnyi/GM6g
cNump5ryjMT1trefgH+vUHg/5yzpQ/Lz5gc/UuWrqYRPRx8pF7hKcgl01qd9l2Pc
gbEbsWHCLz3cSbPNjrg31tOH0uUGa5HzIGoS4HXaw9ChyifxSCo6n/rC/pSIWadw
gXhXoz156cIYRMBsQi8ShI+u9wy0+mg+FpoNnKSw6sdJlm1CgFf0sCBSJffnTnJd
Xt4YwNjLWO/g4Xo7zn0W7Di9BJeH6JZ6tE/Is+BdcJf2x/PoCZWAcReNxlh0OpBJ
egfwbcdzP7wH68oqM/cGf1jI5f8u+lWEmuYPRqffNdq6djuehzSzLtvHXJCnFIlD
74xoXhzgs5kvc8+tbV+LMVbcoTdLoY1VK8mt2TsUYTzICYrx7ZB+auR0fz1zJw/0
t6IdqELrBOT5Gzrpi0+CtgJbOakLbcM1SvdLt8M9TMwbA22Zw21uR7vQ6OydtyEX
DvV3B/mbz/8xCobr9aXGyn+tA02+NuchbTz/pfozrgIXkeTg/0VClb1aMsdE0DYt
c0FXX2rB8RuuOH41csCoYrRbftJI6/haHkE6llK6V0RBxs6Z9lI5tFkXndGQkMti
947FMwuiOaPC3hsS/T9Yjs03Wkpzny1y7IQ+2jW0MBde/+Mul4h0xrEyB6IunOzJ
zz6Lg6wCa6xvOwzClalUJ11kfRZQml+33XVq4OH6hCzcU+tIgkGFpEos27jADObA
gNiBnsmOieaa7HcU7IOCwFjskIv0SdhBqssSclHr4r+Ue2AsM5uJVS595MeaRkjn
05ng9Fj9nKthpTy0UykJS/EN6O2CT2Vn+07WUmMe1y2GBvjsBXvnfccmJEPHr5h0
Ev+NyP6W4neUNbmaJsDRzMRd5mpmvh5BF/gypImjcfB3s8fW+VPm6ZRlVi+v6QvH
aJZWK2HWOivCPtChlsnkwx5DI+5uH1KVgFfvtwCYZFUQcidHYLLlOk9q7zjr+mab
7qvk75qyHRWYocxBQcRxRUI99iZQDJil+KxC5+LMNmA3nhIqIwtCpaiIe7PLhToa
U+PWrfsZhT6soTZVWnwamTolOJ4/rjlgZIo8OFjP0dEChsaDNasQfnQX+b0P/xPC
5kISGDLYXbo78nnK7DlaP2P9WKe4rTat+ptqQ+Zyz6zxnTNnM54W+TWiACETw+yV
hcMI/hGJz1VFvPuq7Mw1KX6m7q6C+os1+tzWoSMLnUAu8wYztfrJ+p7jIeJjZUwi
4Ndq4KQUCZtPWNzRwt3uTmiPwsOAoTKaRMitNsncZuuj7mKj7zu6sbIdNBK3Q0Iu
Eg5LQjSOQa4Im3kXfpnRTcO92e+dnVv/NEZM4wiUytVZyzTHqeDPxrqbkrK55zzT
YUm93/OFKyX+ETmSHuH6F0Me2CyqaLW8Aj7R1r29F6CUTYcFhnfaA5fgrddafG4i
sQDKogvpuU5a30FveYPyy29FZiUL4xlQdABpRd7xFpLqVi0aRQ4Fd+Sjc1IMTdPp
5oShVsOWoyLQziIcduFJUVlz6LMcVW4VKHfyj7ZSzvkoWvw/I6Hbn5dpKhtCI1wg
HKDyJmQccFCB9tzq/EEdzjxOsJe5HsfKGIGSFUlJC8zrGrKLfYviCdunLK6plOYF
Q4FYW2Gd6+J5cCSE8eClHbVXiTmuUyKkKI+E/PNYuiSJN++6NU8WmKgJwdPQ6YvL
fp9pKdlAIP39ShOLGdantf670BWQ7AFig1pUddo1Bpnpn66IyprwVp1tg48AfBj/
2pG9/3ApCVcEFgr4Xrn7VkyCzT2cx6U+HsEacFHj8ZYqKcNjMbsMHIAIf/CeTCLf
nJURbYH8ugze7rmPUGxpE1xltJJbBvUodoLOgPoNcQy6x1BUjZ7Nig30veazCG1W
vZDlJ0lJMGMYcm+frjmj9ycSo/D9wFT+Oe7azZWvIDHDunToJ7VBl+RimhqhjVMk
+a4N42u4q4CalRV41ODBF7a9i3eZBaiOUXA1uoXbAWE2xpgH2WdVXoPc5yBMu4Zp
BjlB7hUpL4e4M3UniQn9QnxnERD9NNBE/oe/8HEp4TiHoGvetImCkHhateDinPuN
Cer2SrWNBqPmv3iwqn9KgcYRdLjdVfs+snc5pUx3y5VqaIIbqHVc9tMbQB1ZLMfP
JXd2QEE2Irq/K6MLTf6CHUV05RGY5RLVxVttf6JRhzWWMY6h2YA7zQWjmZ/mZgKg
DqA1bGq4IrdqcBxxj5JUyQGtyNjRYlOSdLke1gvhPASqpivlCOh9jl14BsCOw8RS
UM+nSfSu5zneYwH1J6UO4Fi4ZkAZZWs1i9dVVhsgYsz2eFdv46XTAWuw4stDQyuc
+8DWK0neW6gUNtghxJk7u+dZhuCK/MnQHFiYhkfucn0TUud3IqSqLqg6A1CvpUnH
E0F+LxyUJrwY+0G+i5Yaws+8X0ITrAKBsfe7NYll/Xpyw8cRAXNogm3lKp6rWI+t
esFNdUyrxuNiOAFbI8j6YqHxp+FPaN8fvBs4EKStWtOIirYfII3RLDYgXPBwoEcm
p8qLaXynaaSnCb/fV9Rf2V25f8i6SoWR8mhUnCeWnlxe7AscpgZQ+VRGnL/4QrBn
bbpl3nafSY6lqFQEmsCkJSCT7VIdpEr/Dl5A/0brGZzLhncC2fDNHx9du7zwPd6X
94jE8nAOdA5Dj1VGMaxNzxGQ4ZFOLYIC+VuPd2ElvIC7YMuP3OHDfyUf2cOkvcV1
QQIf0kHVjjF6dNNVBrNmr4IeasToND2ij/04ek4BuWjB4P9olfrEQMR1urzO+3Oc
HxoXkjeoHFDXbncoN27XiIYdxHcnIo52Cfev/RrbaJN6icxsVkO8IhjnPMv9oIpK
euxCVgYYpdptvjzM2c5rKI26V8HV7TXV4NzXSgibAcxmAUzd4ZE9jTZybdVbW8pk
6mkw75S4YSJAZWrqReteVcSONNf3wVeakTtW6oL7y1T84dF+j+1dV+OlNLBk2ZBt
skHUfHYQhoz9pEohS0zZGunnymmZ627dCM+R04H4R9u5O//B/mLBOuTTzJUzuPNw
03d9snhM3v1/UM3V+HyQsKwkFPq6FDfXTMX2NLjaKgV2Pjsi2lEQAgG7FwlBURpr
fUG04Bxv7M8xCnH9VluK26N8FOND3+DgGopmiFEZj9Smzhj98psQZtVghsgI0W5t
OP1fWhVNhPmtI9D3Qv/PblvVSGx6mZ6C5MxXS8ksBKWalCqOaxXD17YT/7DRBFca
6rNgXatdEb+r9F/kgYFBPw2Df1j5r1bLnN+pPsi3F242pkyBaLUu3BdT0ZW+8blS
FbloBGWk2MgckRyjocnMub+r8dRH59E0rW8XbtxKfjPFoDJ+HEnvd05ptTD5KJvg
JeaqWF0Gg1tw+XzinoRqFA8EykljfceY+bN69FhQdYRWkHTTP+CGx0vnr+sukcpl
mE+hO5ihG3zGhDHkefVfCyg/0/OkxFzY1YMgRzxT0TxOtUX/RTMtty02zrE0NPR6
5Il0z3VqDMH9G5XXSmzhmcNUo9Sqjlpzjnq9uJL2Kf+VgUBJEcw298XZCOYAP1FN
NkITpY9SUzn/edA6O9CWe7yTzMduIEBmKFPvAUbHt3kcdjQZ0RIkUwOTgP0lMgYn
dMJw+krRmvIKR3pJbnFmLOf4VDThaDM7dSfFXtagfpCUqTL3ANxe1Nw8yyWomMfB
WRmKZbMSbiLfpCFIHbUm23q56AAfPyoG9rwFpnCrlsUCW1Raf5h8UQPkeIxfB5Cs
Q98Zx1BaRvKjFCHjQDu8Tl/VrxN4DmHl5K3c/yqK16Hz0wOa9RFItdK0yQouEcf9
XinTRK+6FlIm8kO3M7PW5QEICk2TUsEZ7CKq6gB1vtp+2Fl7oX273/1bR9mHWhhE
`pragma protect end_protected

`endif // `ifndef _VF_REG_SV_


