//----------------------------------------------------------------------
/**
 * @file vf_q_typed.sv
 * @brief Defines VF data queue typed class.
 */
/*
 * Copyright (C) 2009-2010 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_Q_TYPED_SV_
`define _VF_Q_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
RmWUhUzP6Jl0w//TKsJsNBCKqtw1JDv59Ncd1DYtgdGaErNRy2SP4B0klD2dqlEk
YN5n+Vh0lzxJyasKWtokHuUJdTVcg1QZr9DqRZL8GUrg+5J+vovzfP2LF/ljacK5
NjG07DgT3W0/Uj8SgPXpCBUppkMtbr1NkFNu/L/ZXSdEFoSsWw9qrcEx8TUngW69
RHfxZ4puqZnkmtsp/Tf5kjC/Q6YOkD0PNrw6trxF7bMX+xzc+oI2MWEnKLMe32aE
6HNqe+M8THrI2I4Wu1T2BTn1NjlkDurti4bEIDPzZViEwjjHEgPatrJrHKbFSSsb
sd79JTl9SUPrlBxRPfrzdg==
`pragma protect data_block
pq0YF7Jk6VpIhsaRPZuoSn5f7LKMCnBiH4jg+gMFrGRQzORcmWnSvEme3Csvo8ny
WqYljSpVXQoZpRHXf3hM5UWtD6bEiHxHTYDWTN5Bm4H6Ot9S+GD5UZd84wg6J6AS
Waia6Q2Y3+YuiIeRzRZvo5VvJZzfYMn2vWQyvaf+BM8aPCACmQ5cgZAibRJTAc22
lNZ/hJdqGvZtk8elfeYqN+hbjQB5UXwcbLI1h60h3/j0tRf4oSSp79Ikiq0fdTMD
me7rhMXKl/YUCvLdDHR7jGTxMVEQFLh0DQYIWM/Aqwf6zEU3TFy4fEIZdP0eQMlg
fna7Vq5urQbx628Eb6DYVXTjJeSckbaDblKhBZW3CBonhw4M4TUWMvvZjRZHrJ08
mvdHXXO094yBQIzQa4ulNdeAzhlhPEVK8Rkyu3DCZatoQQCygcM+fDIaX6XHvjJG
54pYtUpBdybNxkmHurt3Vr6pxbL0woU5SJAuwMJ+azUmMUkLLyVW+nlcvjE/5eOo
3wyxfDyYqWccExeEW3uBe2LCuQCesGNJ/ll5R3YLyEHRJl6TsNF3DhPj6QLHJOYr
DBKuDglVXjhbVHpewn8dOnOxEzYs/Vg7jjwN5ZbojxrcJJvDU3jk8F8F6pIdfSNk
Le5U/YDVrEPyDicT4KYZpvMx7xZfsNovvC5KxBdAACHfmFL+y6cz6uhbOVN7xKwP
5DexfjdpKlmeEfFbFaA3k4wL6rfb5USsSH7icZIOmOkem6JPqv4q/iKm0lY1TsDU
DAwG2J8Al7GyhIz9Fenyp0021rHJ+gtO9QuaLgYTQDsih/gTgFf1gbxVqh6mOaNd
j8EgafdOcYUqYWDPU9msZWbN2ffjvDjpT6YZK4gTE/BvKK4Av5/hUxmlnoS+1Szm
YdWxfRZjSx4G40usJx/kMGIQuL3Qf8C5STRgiWU4v7LwHexuuj5aKR0TcFrikVHi
tV119GbM8IkQ0VGP74KGaVQ4YdPxaKlHAVYUsrTJ4JFfSo+3X5xzYWl+c1Mumygu
T4mLAitfs02c+QDeAINHli0Kf814yEnKgdceWVZqJmzWHNdSnhm31Q7ed01mLTr2
NEYbuxzjbRGAWa5swYFRdEzOUs74DgrGPnNStCsBqwTOkNPye78Jxs9DdBNnkOhZ
mJ7b9yW3X8bxJ/Ljb5Zl6jv2SVnmsVTv/cU0tCSCTQLz7Gf2NOHF9sb3uJHN4CfP
W6wiBkPzsOr/QEwdW+9rnr5R/nijcyt6gjFedUB1TAp/seet3qvZlWYHjOr5kgh8
ufinstm7TGFciV3EoRcxQJpa9ww9+y4mt+0JhtLLBOOsPi3ZnTrukX9+OqeLhxqq
FQvNR2TkEeNOQ52/uQufAUU6mxDvihqZ8O8xDUGbS5tG3lO2njX2ztMCt+a074kQ
NFCxFdW4xX/ggQPPi9WxaiumYmgEWe/BEncsLDJGZBVvUf/o5w4R1DdkyeVpo8kD
nR6+F75f/GFxT9Kf9KoMXKav79nip3YXEh9lMMMx2n60r4uILaBnBIeMySAK3c1l
haxP+o9VJB16TBspaMCHZ/s7ckVdMEh2r3BgbYFsaShRoljflU6dKXmOI4WtAaeY
0vG+vvzvUqDcpJp5zmmMuLPV0mvj5M4XB6t2emQK+aXmTS2e1ExqLUF4iUyw5bia
gYoQuWbSJAB/Uie3wcp4xdV8dSfR2Rw2bdtjuHkCquPwra6ljiwe0qtQ8j4PE9fS
N2WGxBR/i9v125AmEk03jznaWObfNk3L917PH2AS/6ifhvI7D3Nvg88ePvh7lr4B
6TxIG39DBNDgecseDg7iYfT1EEmJJOE6IlHD5ZbzDQcDwfNBaahGdgeFonGrMSzO
WJnXPr+DGKx57oVjSuE66+6fuPSdzNHFQmH/RhtqkDcvX4pqXd0QpXDjbaaXJI5g
gzOKV6s5JA7ThVj3CrhP0HA3z5eMUrL55zGlVW4CH2SM/TlfgzZ43YBr0+n9b9P8
jSvZLawIujYAbIp3VMekt2Lz0qK1990ytnMQ/vbJZaayuHIk+kPPZn9mCBpYFeH0
EaYs9cPn5csjzt12ikFXmxZPyrg6BPTA6GxRb9P+gzsc66RhgSXpXJsxHT9Lbai7
sJlRyNwAfHdYrmZnpomqXJ+fJOlho8Ed171v+A4WKVSl/A1opr+NPnhK5u2TMHHy
5A3l5RJKLksE6EOe38MO2XIBBRaZF6crv3qoAY71SN4oO8sp60aCRPGzvB+6/kj9
PFws0wqZ4d3sN+C59/EDcIeK03jy9ZYs/ujNbjdAAyXL3mk2sMvHgUEuLNGTIrvT
alqkDkxv8VSil189NCDUlW7Q6jG3qJIpwIPByOQK62qsRxrZWwOI0ViXYTYl+Z3Y
5Dzt5kSuNCMXr1V2JuiDkbjjwksg9PBD1lkQ+EKXF9QxKIBtqq8SO86eANe/5UPa
VucsyHV0RpnTyQ3FQ0zT1cfJyP1IYYA3HWRGviQcvIajAq/y9mPologVW/NH4zmA
aaGAJCYXeHDvCalK8orM5MLIkf6eK/O0cqytY0dzTfXVXuwDWnNb5WOTV5RmPxbM
zSzbc9XKJYWMMs3sxapjmW3+VyLVK8gTM4bpZzCprI4eXPFEKRXaDBZuuZ0AoawE
FdR0br8Tlnodsb2esbjDLMdnwlXIKE6BgEip6bh2PIyMz+flHxfSbECYr+hxKeh5
hPxv7qS56O0M3D6dk8CzzFDZzTq0yUr3IB8vhxNH9lY9/bimezdAuYijG+SkvKva
0MoDNbysVpX9dsXYC/2anQhSwC0CcegwBWars4UbFkrx76CpP2u56EqmJIdE1Y2V
Oioh2TReax/oaiAN8Tx5UST81j8fYD2T7E6iBRROgzpBA43Fyx5/WX73wlXrz8xO
rl1R0TPhfEBB5LWAiBF4yH4cu4YFDqv1SiCViaMvPIlL8YF7LqDZ6VNvZwE16faT
B/mX+6WR9YRcgzmTePGvglAC+VcjB2GK5h3OW5+ZJN431EYjrt9mu1fQTXxxeIKC
xnWcaebmv67NoASNpdJ7Stn/hWOdCPQeoHdW0ZbBnQ7bplwjPUMUOC8xw7ogiNC7
RLoCpcQQXwfUDrXLK7RtI7Fl/01wnJ8fhmbbQW4htn/lg1DNkzi0/ynmurlYNFo4
7zdnj50zufn2BcgKaA7ZZ3uBsujY9T38CFImsmPXjGyvJcm+IpcPNIazHO8OojlF
hyU81u4H6fOr3LGnVdEoYP1IqDJcH9HXNoBLroe6zAZK6uVf/4mr3RRGMJ3v5cWh
LewX1DN+YUjbtNJeWgqy5o21ucYihbbRivklucef7qbIrbwv54snZrbeaSgl5SZX
KSbMP9NSYcXm3Tr06p2v7yNRGrKvvvqldvK3BWrxqb0NAotLKThMt37TchsLeM9m
OBM5YcEo0X2mcw2a4W1XNJEce1GGRvkry+olhrUcVwqCaOH/evaM/1/0aBEdktri
nW1Lc5rSHx1oaafYD/GCMnwI3h1XrS9WKbwHV/dECiciVqUSGDYa3TG3x/C4XnJc
qGe2L4Bm5WKjuVPvh7CYggQAGiNpwWSkWuvyfOLA3ad/mllgY/oymNTMJ4NK2fXY
X3s4qOzqrpdf8MihMtgXqqhELj7zmsuh17AhZtiUprGZQ15cOHMAv8wFFrJYyyZI
H2WXUppjaVpwZpVQmIvjOx0cdP8a5iTNkSAF/WWNsc7dx2KL+dtUvIjCffT4z73B
VrpWDrvjOWN/OhGkZomsdS/BJa5E+bUElDz4tpGx/OHWJ1X/8+8/dYvgGX6QL5dl
9uBd2YENN4s7dnbOibmfysm0wnOh4Ywl++XqJPIeEVh37N+FoOkgUpD/RvjWbpmF
16rKcumFA2PwpUU00/ZmJ69G/J87YnZNKoMPau+OJnY8ns1Jw5gbs07jTp/Ey/Zc
QRY06JSh6SLf5HM5J1M4d8VwXnTaOjwPqsoJzprHr7z6Lhch+ubl0lUx/ADH/c56
lWDg3QtgDBzOGEN6k5Y9IAslZf9LI5xMsodJg5X9iaDrgEVCVElwQ96C8fVno5B3
sQ8UFRc/PaouHlgvWQZmMeAqRmgrR/SdYJAT3r2tUw0lLt20hjJSXd7PcXS1PKAZ
NgjOY5LypDCRLVWAnvpdY3/lg4kriIRXqXtUa5i9oaipzt2kpJ7EcIHHLIH+Czjf
AcrP2QgDApkDjSYd8NRsu1D6fdI0Qvj0iBR6poN3avkMb7u4hZ3zTbj49VYIy/gW
qz1zRFYWZwdlQ65RbHy/qgVkNu8mQLe0lr3Gu+Y7iJEV2//XbfxjOEleodtJ+Fn3
LyKPy8dsIMTdSRTb3tCXRLxr76ok7LUkpA8QebrMFSuGZCsS/QQTZKp+OIUUVxHU
ZGNtbFXaYs64tC81/OCLazProy8R+yhni7O5v3YF7e1GEXfkpYgZFV5zXbndiquN
7OUYn6D3n28iDGXbZ9c5VSYZ3OdAxuCPF9EEkKaEup4zh7juEgNBNF5yxLvvzqEx
vjz6SHlbMLy5+INK4NADZGDexejt4jPqXkRJR75D0p/42ztLX5sBTZFQ/58R827T
eH1mIpcPmp0am9mzt5OrkM0gvpVvTU9rwUOhFErXqiMdObCOJ651WcFxQ7fYeyfB
WU3/aHsAJ7+r4lQTgjkzqSQcZXhRWuyW25KtBiZCmzIlJaclovg2Rr6RYipX3MbR
XkwTaR6QPpqaqwWuTf9Q7S+VDGKNTjMOpPvssxpCPV6n7o71y8cjV14SLXT+IGyb
z5KCtCKkhGtqCF7Um93Cah/4aTV0yFDNXeKjom/XZ4di/8ahkLJDZpn7gOuOjDDV
LRmqq/Nh93/MqJ+D4C4FlOlO3u6gAFIVdNmN4WlunG/GDaF5J47TAQ3eViB8qWUW
+YXEbOHQQAIAdyaBSO4wk/EBeYu3PD7vPVk0rMIEyu9uA6GGFChjKfH7Uby6tj9G
frbNfWK4ogL78abskUy2ScpCxOF+WYGzX/qtV7UxlBoNUTMcuQui0bM5bbVv0T83
WG5YMgLLbFjNY7gvtRR2shIUvzRMrMaV9uBjAU/otWon/CErXoataqFIeHWdR6q4
En1iedvlG/suMSSSl7Nszlp1J4zIowleYrwJPEScJf6Nzejhb+nCT6bbtfvMfvWI
XwMwy/Dx6CYHqM2Qu7/ud5yQEDWcKsBhEWT9JAaI9gEDBiQBTgKFmGuJg5CmN58+
cGOBIDPxefQNORpCx4ULa3URI8aX48AzvXmU3gD57HKHKO5tkXkIxLJFZjy3C8cc
xGa9faQ+cm1DzDEDoEwjcHG3MX2k4/SlZpwu8fhI46nhhpV0P8l7ml0eoIP744Tl
gxxj1WFRu5sfOKzgOsvomq+hZpQ2aOxNaHcNPOs8yA2f5OxQkcqXHZMg7ieJhMIB
I3tuSkcEZ28wuHEaFx5HKeUBgSSXT2PMvzFPrGbmOsc7tu3MuT/Jg08vq9T7BCVx
abKWOOATuEXvZbMoG5hO9df8zuaC7ohisoMGzjvVpfVBuLW93Q290zUBn4Yi2YhI
u1rVxOnn4+QJcVmtNl5ycmDa0Dvlax8cfYWeSXQ6InyWmnyMsZ5hexADOetlD9Hr
CS4/lB9KLLfrVMSUuNxpO3WREQg8O4EX1XsN5/p1/5mzHMjTpWcHMt0Hq8VKrQ9A
0aykEGUjdIEZIMxY2A8ZNroDliKo3QZ3IY12slGdO5pmVpmmHvu3+5HC2aDm4oyq
gESecRd2R2rD45NktEMYclmBxasjzlUTlmI3sYuScSFdwT91/WSgs1epuOSzSbWH
dwdIsO8rfAIfZqtHxHP+4GAANM++ZA5Dx8LU6XbLf5iUNbFQsgsUJ0TkTD53nyoN
HCKmEKTFBJu9L96vHhZSR7+5QJ2VuyTxgihWc7Mkj//CX+jqcq/qQu5hJe/PoEdF
M7YxymIbcvCfDN2mOaHXB0jwJmcgHnPD7EpEsgiq78b+nrGWYxFxVPPGw42tBBU/
VaoGde+0OkAyIsPk68epaVKRUCPSUY6ObAM454eseEbx+EwYjdxL8ylKbBS4Kc0h
GhkS7hr7gRsqNrScGSlq7I523PBZ5jiw6P9gfZBFVSS15P/cLVQxKoBxT2GjN0e1
knoztYPZY/Yu1RZjx5kUA05q1d4yXkzMta21WTf7p7xGg1ZcMkWPbIZxhUW+/6hV
Z+KktybnX7hVrYecmvEvj6P0dteT3NRf1kPNDT7jPDl/N20C4dz73eqSzYOmd1p4
VJt969ZOX/IR0Iqqgds3Oj2e5HciuuxBf0SKPYoVFhs=
`pragma protect end_protected

`endif // `ifndef _VF_Q_TYPED_SV_


