//----------------------------------------------------------------------
/**
 * @file vf_addr_elect.sv
 * @brief Defines VF address range election class.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_ADDR_ELECT_SV_
`define _VF_ADDR_ELECT_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
DUVE314iT48+MVHFSd/ZfkgfS6yHCL+QYAnjaeIO5g96n5GgsXzIQMJc1n0eqAzv
JYuxVXWePaU+RJpGMFIvC8wjsbZOusMcZxmJipi2MKP0kPwcaE7c5ZMewT4+OE7M
CqpyTSJMGyPmIOCmHk2aYEkjN61T1cv7QsqFL0+cEMeI4XnMugXWqrQjJ806d3i9
7A4trR5FjqL9oFxmdN56pFZtkrvELzcTuOr1+31P5crWTwi0yIgZ+LhPAbn3cIcD
7R8rA4YzPU0j0uH5HrMOF9Axu0moQi0pPk3j1DHCjRBNbO9nj1+LCW7+v/lPtgTm
MYbBpmGOSzaIBXv2wgtcCg==
`pragma protect data_block
0PkDiCoaxXicOfeP/omrumSU31q1w43zQALYEAEtYfnJleIg+4yCGxXhkQr5iVN1
GJQ7wenGkeMHCy7jbSQHSuayJJdg1VHhc8pfsIrEhzOV56+wS6XRINwSBwqBafou
Ds0LBjFpdeVKjed+2c4vrvXAd7PQQG0L1CwS138Ehu1Su8sEDeSaCcqoZnJpcT6r
ae0QjY3mjt9ozvnYfND0yi2x631EFlSqyLSbN/gXkhFjw8RzhjgfwwKhqraDwKwR
nYcI9329T9vN+uydiZgrv7B9x7GSWIdh129hlUjasgngvia584/l1H88LUg2je3l
Amc9sTzJmu65+ofl9au7ZAgaNaj05qjx+H7JL6RKHi17BVcL9To7ZOEAjHC6kFaG
LhYbvUl9XL7fMUZqO1ZcRsfs1ul5UbkMFUPTHmY2ue5E6LTOI+PFSgVxbyAORdxW
w2EgsdA8l1BU9YV2/jyDPthm+9h+MWnVx0Jy/jmx3tNMyAoAJdagbtLQDXC4wPWo
BAhjGJuTN2gcp/nu745Mo7wAnLCdra4sre+WiBuHB239zbfnDB2HnvFFCRAHNAEE
vNMt/JX9tebvDZ2OOjHjAo1VGv3pT+Xikx4Bwrw1p+Cguyv7UKtnwoKO1RU28XVf
PYYtH1UP0BbsLBU22VcBroZHVPfTMPDb+ecBn6DiOjRbWVULjmNHh2hyO2SBkGdH
YiSja8QbSd2FzvrUxtn/N5TUmGPWN2ZYjoKXss+39RY41UlBFyJjlpcB06IjddKV
gM5uCC4dsCviE9yG70/NDS1iqAXCVxdhfUxXwD/N0TEIcVu3o0qURVrUqJFOCzBo
jA/hPCpb1IyxE+ALo2XYOuRXiGHPPR/mL3jjE3KT9J/nCK9H7QF7RBvoy/YONnyr
IIZpHsP4xDzrLcvFf3E/8ArREx1KHgIwFu3Xs++UBcHYxY43QEVNkejaZkIfISfY
s4Go20BTWXpcvHFPMpdWOXS1LpLdsIKm4w/GBtYcrjnhyf1FuhGNLdtN+xoUTtyT
Xieo5hlJix0n/7DftkCS55pUM4PsEP68Wu3vfIFlv5t6nlfQYwu6zEZuThT0LNVv
+XXov4wo4yMm9fVBnQf8hDOf9HedrERjT0FaJttVMgOdH0OJkeS/fUlkoFBLi7P0
z311izXS9HXUGkE/lqvv8q9s16xBeS9eYGjT0EP4gAgK3Vz+Vz8vbzFmZwnXAJai
CRykAphrrUGbzrPILBLopPMr7fF3YhHfWpbqHdMIT+ckyP0ETveCI8Mc/Cd1fKFt
7A12tS2DTcmB7UXPzCWmrQiS+H6u0KKV6gp3pJPiIfdyGxx74uFcCgU8Qkv2PNHs
mF0+nsFC4FbuKtWdOoHdhRaKOnof+8AyEVsa+e1L5Ou6pfyk3nztJRAPpALEi+tG
5KblNY99NhkBkr1ApqpvJiS2b3UG8VNg6VEgxvOKBe3TrXqMPWCyAY+cC8DE8Gyp
Sj3fnlcR6Rp61oVVKHV5NLz2tSCAHzCIZNvzLthWliTkGQdsDrzR4WCI76AmCZ1V
HktG5RLdTtFtVShOUBX8XR+0qquNOUZjaDZ+/f5R/khFC3C8Ri8msQr77eOD7H5k
hYzey0WWjGzWnJASEdMiddf+V91BK1u5Pk6TyF9Mk39ki9uHrImPG9gzxYeW42+F
m68AJnLlEpBjU4ja/ykluA8qkAjopLQXb1SIBIC372amj2u+5E2k2E9dnL+nFzVE
uS3psFzM4oneUqutECPNqwF+L/l8jozLeb4BwGy+K+7IkDh2YCgz0pw85GkN5+E0
rXVWdbSRZeY70yhVV5HYH0ZhTbuvER6WYaJh3A5C6f4gPFNUWCLAVgviJkftwtg1
Wsgwz4oJn2VU1y+Typp8F0fqUWDBFhIg08+LhiFUn+YAiJ6VwUnYZWNZFKmzQVbU
DCh0km9PiqF/KPW4pXrStaMhXviArkXGKi6tfA3bglQ9i+WXcRrAS4uwjUYWjW2m
OkQpcGHEyRTJK8c4Zm87iaNLsd38cVVqFmXxp4gh2ngNiCXUSOLuR0FtEnmSePmq
zr8GCD4cpyscOhE+keki+1O4zqj2UwOPe2XRb8ANUSj+Zlps4mqNv7QHNuB8U5Bg
XK3K6CAbtxgrTnIAaK/kO2k9Xt2wvX9RUJYeCapg3JY2N/2xHW4zNp9iN/O6RXQ9
BIli02muWVotcyPxf6ioNqjlqXNJbDS8Q/IKmeE9Cl/ba3acynFzUKQzJ11kaaUD
FSKfQtGZpUd8Ih3u5FDN0nevqjY6GApu2tOXzOSDRl8ZLK7Wks//HGDWQnrggMmS
XLJnZjpKoalpy7cNjG/V0x3Wu9ggbNLZPgwn7kdqqLwPw6s3Y5+Oa+3YoGI3e8FY
5vcWgDsqS+ZmNUPS1lodgPsKgxp39hVme2NcmIuEyvproHid6isTAEPYbDt2KGca
K3A2v5KD1aGXgWP/+DJvV440cZYUsICaCQ7UGn1NnuCAPtFaLQv2G/Q3mN7ilL87
z1QhiT8W9UTPdwigiCdCzBkmwN6YPjeNfH7pNv3M9o8pUGVoUeOeX2Jyiwy70OAk
JZtgCeOSXoMXYXZXTMZ1J9k0nemQRSL79X8YXIDvp7sSYo9dQJ3PG9nN4dj/pokw
Ko+14TVxGCoAh7KKe8UhUFTi1sL5czYHgnnP11mzJJ+NvMeYd9xqR9UzBnhv7JJE
ozxPFEDU16qw6ihvBze5AJ/Gqear7YWlBe4O7QwnGrTs+UeZEqLitdr+1NkaDjLj
dOicOdOQ7N1FMM09UsQk5M53Iz0akwQ6FTxV9kgloEzQlm8MrIaOaEmacOnT4q3V
1AtZd5W/L6rzUCq4KvoqYzO2SiDK+r3ZGWr0XlFxvfZVPJfUNIh9TkIJL7ccfwBy
0A8s/HHIKLyzamdMXYO1scImvL1gRbDzBxXAHIC+6IacMAZzLYUrLq2mHuxlKb0A
+Tt79+Ja4h4hnYMkMKjeTVAt5aQlEFqti6fQBMNOywTbZgcYSsTRI9mo7Zw4xhIZ
//j6Ug06K8nnbGPDtuEN3jEgj1ebFw2nryQm4SBhoOBbYxT2ftDRvDKySdyp4Txq
KfKHCb/mJ/Ml12M/SoCnoXNLZQycLvdgZxYDevuzEw2L7eZP2/wRaBRRUGIrwcWW
RXzela/GJVeiRO72ncdqfkpvt2bWXccAv/hhY/inc9wdgmYy/msCr0Z01B2w1t0F
YJ2potInqq05rBiHh1N+WBkagnghMGXonZwfVQzSDjkFqHv0EBQ28obgb3VbCoVR
sDoas2vqGfYPhc2GD5mJwYMt0msMFlTSdPifv+BBD8iXI/zfHdWPkYbirmDkyKKn
fw0FnuQ32HQoHqx7rarnSOcp1o1fN4a6CWG+nWgJ1DU4+semaDkmK5jLf6fMDRKq
geCBirF1XDKbdQ3x/Ml+X9nq+uCgLt6+JVWS1GbDGn044+4D9z+wfGvCO8TyXDOh
7LejpCy4WOUhKpKFqfhn4DaCnRdQImqC+xiU5LA5+d9yz5JEVHBryKPjrRxnItKM
MhnmReDtY4/YHBw1SBfZ2GyjRHo/e+ehf5KRiRXklc6XUdOyu/SyolyBQM4LAMhT
NjoodyxblXrRaubYOncMJZDDji+DK4AiKU44pVqVdZ5Ens7RSUByEBEYVn8SvlWK
Kq2Z+nOurpCBJliKyeM/63AbLz4jYW8FErdUsIpCHJNcsbBLq7h3bUOh1n5jek4Y
Br2FJqNr1arKnx16rDUafkunZUxO0d21flFglxL3dx1kXd1ApmKKB4OsOwSFPj2s
SuWL80l1gPnW0efcKcabnOL4IRjEL94GjDoh96UTQ+jdU/mu1EeQREEU6L9DY9Yb
mEsZZU6kNk/pF4paTdSg/L1tiUTv16SG+WpcKXRoEA5k/ANhxh/BYI789qCCJaAb
Xr57qmObv7GwH+h5aKRNDI45mXk5mCmd+kfrH6Z6mQL+fh2OH3ejX7WSS3dc120s
EFZRe4sDl4Jeb/9zZqmsHdP4/ze3o7NUaR98oZk0ag495pcLMxqZFUrQ8BlKrNEX
gnwU+zehWW+0YK0e1eV/0uWlx6nYDHOM4OcpMvD+IoFUQN6AwIRrvzG7lkDK7h9O
dwS4N+MNDJd7L7NfhdsKjsSdfUDsHOs0UqaSVH26DfJRK49eok9KCs9TpLovXaOC
sE0bv0ihKHw+praz20L6xnsihGkQ+G0QK4V1GDg/pKeUUhigvf+L+fM6XXJHOnGD
q2bfJekvUNKqPJ/NEHS/2iCKhBFyiqpCLQfsqlpyIFPBkFoXQntCeiIMElzGCYBW
o8dU/oCNMAh5S/SJLnlWCqTRakiRbxZxT/RACmhetDh4XCx6GVaqosPPf22tEmeh
Gl1jDdB9MCra++hGsCkj3reYriqfyKS11oEJqZ6oiKNchD6CvJw46appRMqaEVuT
wSX83FaXWME6UPi5L14slQPK03dDvptjq2u1DBV78WpifP4OslE0CzY/dMbJZ86r
4OjrbXoOtLRqJrC5m/bbOiCDbzzZ7D/MPkUkZaEpBOfObbdNDwWN957SwI+X8HdG
OA+MCnJ187brZtoOSaLV4j7jfCteSpyT8QspUK3IJHriSLDWHxL5wKRMbnpRXFnA
d6OlvxLeFRQa7vwsAB0bAdM8qU/SF/lwSGP/GBUZHEPQjJALbnvIge84AtzDMZwD
GuvBbA0ZWa0Y5s54/9Gaz+sKkhjbEeuLvM/kp/S8IHh7LpG7JLCQcCr47ChrbOQT
Ri9bIo9qUUulYlfxmZwqIig+VnlkddlWHA1LcVbS/CSQWw2jLcFCabPOM7CD+Z5O
JZjA4m2qmLD46xb5+hUwiVwi8XbI3bgzODtMZsYnAGn3DJ0VyAMyJdyVh+fu8OA5
7Ea8dLcAWcFIXFeszWYF8gmcYmFG8GdW86VXiAR6gQJn3egJy9TZwqpMiwV2DVrX
gUcf9zSUt1YM9kA8rjH1Q80WhF2eqkhlKqiN5BPK4kNLoTCeSjvqHlk4uvDU2749
nl1mXmJ4pvsC2EX7+IMmyQTfW1bcIR+YkikUPMnvYC5rOr1LT+35MSpjxyNoLIvy
Tce+5XzY8czzS7sxgukNMj3SgZbdBl4C9F6F4a2KZGHKHnArRXMCN1ck7hhJVOgF
owLGr4MO+f28ueIoSABRLie0tql8W0xVfP6qNhYKpkQEjbGHAa8wq9vZKZHTbtEs
K6Pyck+Ss0gF9rnWo6G7xk+tkoIukLj3Sse0N2KpV0KKRRqL47DQFkhOzWDS5Pei
K7Hb8WNqrr09HLalXGEMvq+hue/F3OQDHp4fnVmxlzAr20KuKFlHVaAtFOcvUrQl
BK2ZHYK0Udl2HfcvKDwOvXPq02RLmR2sZJra+M0tEiCVKSghZdmXex+ep6iyPvD4
IWgGm6UGKymNomxf+uma9h+NUbKpHLfrLiLbGkWbB0YQGc2g5ECJ/F5QyLk+OmDh
mV6DNTi4h2mxc6Vzp6wkbSs7kNKGZLncqABiq9aj8h9tcVzZ/SiPLEBJvimIkq9M
0XVLiRHWwqdqO/6fZF7VbRh4FGy1/aVsnrpDfR/Lekv2CrlELXSGxLavXcwQDERh
geCZPfT2sKHFzf8/7E7duPnhFZ42E2g05RpFnvJnBk6T+z20/nEwX3WWwI8oZWJw
3Rp5dIVvRrl1mCy1WQEZqs2RGJxzIMtHhN2AAE0omkk3ibkVEVLNUhpjnNNSdo4U
LfwNrQOLqWF7lMq3QubM2WlLX2445PYnNqgSEjB7q4F7U6PLG714Skr9ush497I3
dQ29/sHoAFYrD/6fqByj43kIP6Ia0RpXMb7n7ZHEKgXVRsDyKNLoDBD+zdlK/0ic
hV5jNwoHgMTqwK7xguQgMWmbqGjF3Kwrhdmeip2uO9lUztAXScgvyH5wv434ILkA
iitjIC4IAMh4Quk41gn8aiZyH7i7Lkrn/cYMlF0T4wCYEaS/Wqg2wUw5WX2zn7GA
P2uJglHP2YM5eKCP+zLEQE3G28WvHAwvSxjJllyLXbvB4POKlAtXtOAvB0cKSzf9
6CvuY/hSxSynzcCF0xN4H+3zPH2JOwanOCvmKsMHtzSo3kXro98N2GsrtvOwdQNE
9KDzKKn3Zdg0n2cwHM+/X5YbOAV5IxslV7/lz4HDSd5AYNh1/+iZ8il+9o+c5Vu/
Uv0EndRVmvHJhGCLoYqIWjjlUKZkNRLukVGdLyTkdO6kDcLsR7e1+AhbTa/4tIZH
fmmGOEPbepJG7Y5r5sLVCj1KKpXNPiH2k9+QELek1sZM6yzbRciDv85xM27lehy6
z++zzErK06FhOnuzNIBqSr4xibVAGvC2Tzt7DSVJL9lK1KTxgdJgsTU8E6nI6DkE
6j4FVGZvj/qoAizD4NJfyQOJbL+Ahnb3jECdCEfm8IZP7tocrtD8Xyxoqx6FX016
CIBPGLEkG4JeK4pesAiDtgamSYqv27bZaJfXD+mJqXigXKKJAwLtHQNP5hWw+hAE
AABc10zQgcdBHDUlwQW1HRZqlrv5oBOVbnomhVkrOl9uKRHhmrxTy09eFMFq17dC
PfSbcnU6AuxKJC2KrhZ3U6Cd1W15tEwbsXo4bXvFiIAYCry96vgE7/42EZAx+8sn
HXRBvvueKgVVEt6hlIgLRHaq4IVEFlXQas5IL7WKzNJ92kALgIy7tYoZc1+MS+ek
pdmX6p2/UKqvXk63yQYUrBdEquc820V/Wmprp6EkcdJAUd9iHWlfOjpGUqwx2io7
la7a04QOd2Qd7+d9D47AxhsJSiK/uTyVN68VxaHc0mEayVMirduaI1TRxNG+5OVY
wmLFiIwNg6HOgEvsTVMlkuBk8qrEegPqF/6fgdBFBTLT8RHqrn54VJRwhp7C2BOs
e704iPrYdVHB4NKJUR2pqgCgD7WwdHPOsYHzpESnA81PXmNMrfrout387XHTcoKO
MqmcYbRrcHr12TVqLEqkb3Yc5VfpWmPxi16t+EdKUIMY4OmkDdYnfWiF+tk8Kh/P
hS/39syvl/9LLlyzNZ5XnoMsF3wqepa9BR2MR0fS6vwGmCgPxvPpT8NCqg2FXFPJ
OfR9ptXVrZwWkrGv7EkJOP96SEbcNVWeLb/RmvwP+wMcsbshkQdAB0j69VxPDNU9
T2XnsWJywH9999bOwFdCA9GWBfp4l4NNOLOgh+r226YeN90+zKb+q2Ex0nPSrdMv
DP90Kbf+4D0CdQrQxpR9JCbJj6ocN7b3OODE5bOZN3Xh7rbE+oIO2w50xXlm3uHK
HRf4jWSGBaeznOBu0DqlBr3A7Q7ssHkTWt4ghFK8sZNq9CTGEN0vquMknTN+GmhW
yUTYPhIG5L1UxZMUcDmRd9XG4eHS7uMpqpcB+pGxPk7ii9SqGg23rf6dphndY2sY
BRUU0yVUqCBDZV4n+yu5JbPpFfYqmoryAqfzUWEPbDdrUmtuM/0lRgOdlnRILZLF
4Qo6xwuZO2Fz1x+ODzqmc/UjmZmvSY/MycE/0SyKa4jaba5LeKaAkDseX4vylIU8
isNRzveYR8aPeuo0F8p50X2K0PkqoVp5OOpsb80Jk1Vwyuyhq+0JO5BvMc52ssss
qfVK0X2Q73kj6z+M5tWRLgoaCjUJVtlJMyI4z5dCv8c1VLkDAAg0fqF9611+Wf0y
/b0ejLM9z1NwGboxWEf8yqY+C4gHYBVizqtZPKQuuy/0W0hM6BzVBUFwXQu7Rwjr
BmrKYBXT3+URCWF5+dUwU8qQPOTyShALwdgIxg/onZm3Il0VinfcTGHNXfvwaM1k
7XYMnTIzm5q0PAhVfQ7xN9NLWwA6rkEw8XNnVEYNZty3Lmvmy+8hvNCH+/yIZQyI
POVuKqqZhQLYUAPPTXAOGF7GaDb41O6BMbOEcFFY6nsRED8KeOtHNo7uZLz5ufHO
73P8mtx5LRyP7u5u1tuXooGB33p6dmaqys167oocExq7xhDe4RP6hkaLc4N2Qs+P
R1ymtsb/NpbN7HNgL2aomsNjIxrLAQ+S/TCFloMRgFqS62JNb6w7r1oNFwjB/iTT
StZBYfw3C4rRfSFVx/6ZIVY6El0IkchXxyGrm6y8a0cDWh4fnoWmKhnclYaIXcVx
BjsPGe+ReyW1mDuUWzewWU8BHDx+l1TtHZKdTCuvPyOttyPGa9wglDoTDLb8+tQN
66tCGaL4pQ1BQ1BCGaoDdwCKwghi8VXgq0kXu/9lrpFU8LxzyqdRh8pwmNH4lQk/
YSoLGm1Z1GuKunxEc5lZmLq+AYZOInsRSjdpDkftYQYcfr6WYai0eMVEZ5UMRNRG
hRSYRHrkwa+2PLPdh0t6kqRoki+lTUvOhO8BInTyuqkslAkveCzFip9JdPg8ExeB
0+4M+vZ5s7Kh2A1Kz1YEI/2Y7bh2x/Q16H+KUX4N8OI6S4akOPOEn6sgN3FPI54M
N0SMJiDMRmjydxIK+XQTIwor+4V9jCi+aszvYdnA3i7UdF2ziEpJYszdQL+nnnqo
ztKKPxX9aaOl8kI1Wj4WUBT7XobsX00HgtpAwsLt0uWl/ZWFNJUCLaFLNmkbwupa
7qu5hhvxlgr1q0w2RV7NZeOb85o5GEjaH+KcoZ4UslZUwVMKcpMGNcnOdX0oGI/I
eeIEhA/vN4FkZBmK1U2bEmmedR9C+37PxtXBy9SR7KozUBOOsE45WtzdHA8Ia0Yi
ymj2edgLwQYlngscdcJ0vNEqt4YWTxVnozmgQOTjvBNyDnAK8i9DWEGqCIq9mfg2
TGU3SN0Lx7FZK28YpTJubjiZTZX7nkW/7WhCYqRH2TM9RnC/XpXo2U8aFAwTJjji
yQxPOHukgBH/5RW/bxBBOzr5Ii9B7LNtmrFqshx1hVuYof+p/75IRcZEAZ3DMgFS
VL5hVXKrGDnThi/ZiMlXLbX1vKLrfrW7Pa7W3lfBQXUGSdFGK+d+3dquqSWcfiDK
dcjCi8alxagAIM+VAsCZ30UwkFLL6CZSQo6DzsLAKucftzR0dBr5LvQvsvDcidyi
uNCHobqqwcGsnmh2I8F0ttwsGieKwXvFGy7nD1GoNIHKKdZHa3HAAWcY28ZEJ0kq
IABt431kEa1gpE+8V3iev1TKv/bRpUSNZwAX12Kb+jpupxZH2P04aV6pcb+1Yd0c
1hLX0TpZipadms8+Yrm2iSqd0ghneiGiB3RIs1BptK4kxUI7Dz05gRv4DsOOmyYm
si3YQLkqm4DGkM3QvvpuS1CSCCXqRpT6gvEGbLueIL4U/yU6e8VRPxfyHikPiZw6
nzTDVlrsCgEhvv3je6wWYKGmIyLsjxdLkd7PhA+ff/prMIaJFIlWYEmFwo0MApca
HB9Z0qyreb1ICO9vvkRTm6wPYXNbhwMiWZn9JtbwuZ7fmC+F83OKczAYxC+Zi8dR
MIeWpowB54tmqqj71lxstEFHc/ZnyVOC/OeZUzIykd2V5mpGD1tAsp5gXLdWCCvb
N35LKUhb2ctVnggc+CSJjm3wQiSm2ZSUz97A6cko2fWkX5YGJlXdEmYYE0Hc8EbM
llrLwnS4eKkNnzmvzoF5iPiaqk8c8redN8ZPUrYtgVfmuCMaYyotWWWX0s19+tBg
OTxv3AwquiwzxeKcVbeR1WG0zYFmHEj+fxqLwyP5HG89aqGbEiyzzQ9vOSt2odBo
nH1uU1edi77qQfNbUvqHz0Av3vYbS3vScGwHPnrf66H2qFkWGBw7YCzPjzIYfglV
h2DcarLzaq0FYdOInozHsvEZNZFeMwxH0BzJr8lAixbDn3PAjTJBWFe7LEsN1QoF
voxLHDLGvE6wAvqvqvH041p7mSYawmbrraj7wNIhK5F2bST+dJHl+lGkokdO4X9d
d8ODDJR3RDOqaadXyQQjFCQWPz2mzgysCiyff9FZwA7Oa+sqDFUNdp9TCKYtBXpw
aYE15QSsd3333svfshDJmZw8EC4mwVe67440wYRFji/5lc52YPpyHWHCLMsLQLra
ggizjDrzd4YtrT6bEkfTtxqvTeRd87rKtpkeDL0tUf59iOSh3gDgHgEI17Xgi6wt
tbEGh+s4zhUNAjk4soIcfOELGwcblTIP9IvVPzIJn1Eb9bakGIfj7nalzOabu1cd
+zcmfq/Sq7TxGhDWhBEUuDZxLFIQVqgESamzw7BC0fMGtn6mDJXkRF+YktSsHBb0
dKphT4e1jNsrvYAhiCXVgRPZT7mf9v0LL1b9jkH9VAkvAQEnC3NSEBTM4ZW7KoDB
vlvV6J+mU0YA+hjDrstztCc6/tagQlq2D0YTqEVDIQGXpLFs6w1ju5JrITELj/na
ZyKfKX/oOIj6DhuBH96s32+xPvlEPX8wdGQiyxi2kHmbfRCMccQH9JmTDjC+m5o4
YG87AtGf/N17XLp8qEd7ZU7P+xp6emKATwW4eZ+Dsdtg7fzYSijMtvKzvQKV12p0
uawAchdcmKC5vg3DDkKpyyZ3g/v2Aih7RPIcaJXzHR0IwLG8B3antZyflA6bMe1v
7GPhVuI09zh5gG8S/akEMRIqAH+A/FR5eXuZmcR0buLjhxUD6pCld9ygbQCXamBR
nqFHMCTGwUMtGy8YXw1sZJuXRwewuIC9A0JDb3yhJeh2+SG/Sz6d0h/kPHZuxThj
xFSK5lhlXV+tfozt2cBiyQhG25WOFawF/DgfQjgGHBcAoG18CEe3ZyFbI7nTt9tB
BEbie8tzL1pILWHFLGoWKR/VYIcEslMZi17ZxskmZptpoqqVH076H3F9Zlauwgy4
ll7Kb5O1CMBDfD4dAhE0YdrGtFEG27GaoJhcy5YYGzD3tUp4ta45ofTO2i2UxFc/
rWEic7YbCo2+eK1fNkO9CHQF2tslX4Yym2SASoj4F27O5Me2a6DOBmzyecWdCJKS
JrGm04+vRcwMYKXETwrTTb2UHqFjjlJX5fo+8uVv/CSkIJqud2aPsCv01U57G95o
9xrWME26Z2oaFzilLa8mH5V17O6bG0anodjE1f8DQE7/MByj8q0lf75p1ywmlqQt
dr7eriebcbYqFcm4aVwUXV2768eAGnV1wsoQkIQ/4ARV0Ob95AKuOKvLLkmrzgrg
yYSFens2+elKpt71KDuYQAIsqSHQc2ExHYJAOAQ6Czw1r4u9icTZKO0K3CTbiHMB
D11wL4UDWoFC5f2WLzXHq+MzeVx/27vQ5lbnLHxr+oF+NZ5rU/fxcTCScK0bNfl/
3Jb95lFb5L19MS2R50DWkbng743uyhdHSBrcDsfz0gNGypXEOHiGGm3T5GKT0atM
kv5BJONFD8E0+WNUegHvbuFx41DOzhWGWeoz1TnDmxZYWkINk489S5yBqygtBlVy
X0rDsQUzMMMmatqVxqIozLbRFyfK2+gyHNWc75V5tGGScbsOBKDKv/xwpf1Dze1E
TSoiZDkdSKy5bnSDZxABB7jgdoZdR6D0gieoZ/reE8Q38y7AyAVGWtNr31CjBjjW
7mI8GOgkY6HAhRh/pHzJg6m9BkOKuM1jhPkI1lFsQbrhc/v6+I/VDIB4auaI+yFH
VwQadqgVyEKjdmYb8OqTytaV8pROliXq75eLWU9sdb65hELL9yfIKzwmcoxFFvZD
UFPC7apP2RJsrSrcGM7E5bZt61ow3uuZF+k2FV6xpYDq8uDpCYSuucwY/fSrCHlO
zQwE4PQ68VtrUoOaricxpQIdUC2ckWlQHHKnOFsUzhTlS3FSO4KDHEWTKw2flAqB
RR+QHky6VezWvhkPecCeVYQaeN9un0rEoBGn9K94TdvUKdF+7JMxUvtr+YNubC4e
EeaROcgxsQVxNIlBqGaZnsXrQ+HMEjbKB7NjdQgY3lmBDShp7FwQ72+lBuPvsEjd
HrL5F+lbtnvTKcjlEsk/+ZD/0zpaj9kBSYyUQL1O03pnohv8z8Qfp78Wdt5CBzEm
A308fr9DHz0Zo4ViyER+rxFd7Bb90eLCnWHEtykkUsMoE3iyDjw5RjctzOODaoOu
YNLar2mm3sfnnUKZrS5YOpKe07d2r17q/mhjg95Q8up/vJ4WZCAhUf98YvhpE/NL
FwMvG6ZkTwtCJg1RxEa4xaHnUNSbmphHiuko2u5oPmqEiVhItNQnQstWwF+65LIY
m3Ebppcgwlw1LM3SS6vsTSXy3mqKcp3L6BMZx5IKr30EsV7E3PA4kwy0Z2gwBuGt
SR8gTUEV96SFji+n1iD6FVmvHat5S3qdc20vj1Kz7I/gHvp3f+hsqxlPe9zGdvCE
b8nxCWNQoBz/mqCDatfYvbqRAav5rCv5S6fwtvAm7NmU5IvpgtmdCUFNu5BEhfvc
/Nb/4NH4ZJnV+5CmflfBWRoldcHbOiI2enD+OnSD5tUSAw0eAtMiKnjkXuqkXqAj
qLphqUbw7kI3NF6jojZ+4K7VzuhmCZ6YSLteBJpSEy8QAy6ogat6rkDb7iuGShjS
7Vr9GWdwb/gYs+xK553vOadQlu/z5R/dY6bWoakFt5lbrSAUGERspJjiSchN7Qux
fW+gkkBbKlfjS75YUhSiMTTDTUkubAJrHBsDbvg3jc0g9H2H8HABuIqKhle3BNE1
9ZZMtBgkpTPliXwhTYqVIRJqDlPd3vuCX3sXDAtkFY0y3Ab4OtGEz/bkUzuiX/jt
EoJUVyrLDFQusxlRVKOo7d/p5D02aPdVr5TJyF6ghcwX82yYZvTr3hKtO7Z2xpQc
b9Q1af0e3NKowHoeJPw+dK2iEz8s4tjFXRT5l7HmMF4ZFbUP/yPeGvLJjKzTzR/f
NAR3LJqPesM3CEEixvRlcCae6tEHcKPx801BzmxfBIffmUww3MLbnQE/VArjKu2Y
SIN65joNzEBwANJtDecEEscMJnZRl8YI9i8Iq7MTLug3s9Qr+4aX93v0GLoeswf7
ttevls4qoNcKqvrEbAgvpa4oxtdw+msGs/T6814oW6qDklS+Lu+dWNq3qFa26M24
lpHAsC5gYJ6oy1Rhl9nQTi49zQaTaAHe77eCjPxeQfuwsOCGIUqqwinNKuBO6fNp
x4eL6/CawTQzvePY43O5tPtkwzKADnrmYU78gJXLByAQzk0Tl/TnKEMEp5AdXZIR
OWfDaHPsbus9iFInLojDTA==
`pragma protect end_protected

`endif // `ifndef _VF_ADDR_ELECT_SV_


