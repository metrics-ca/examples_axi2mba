//----------------------------------------------------------------------
/**
 * @file vsl_addr_range.sv
 * @brief Defines VSL address range class.
 *
 * This file contains the following VSL address entry related classes.
 * - VSL address range class
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_ADDR_RANGE_SV_
`define _VSL_ADDR_RANGE_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
HqFFWn2vRYqgiBVeWk/gXSXEGC4ZWnKgkx59PtNjHdCZ3CybSWiFpxOwBk6QSzUL
QxT8W0FTgfPLkJLF09vNgBp+aB1ew6UR6SAbeM4OYcJXLbeRHLZbIW27IdDIrhPM
mbk81hCK92/3edqGFkNIypg1FDy80XV/034TjthioPNA3SIHo0nv296ZtvahLQvB
9k9x/1NklvM7jefxWAEQN0VPy7aHmARzqdc/Su3KJGfB4TT17oIxcyZmdx9NcG8V
/34YxghOuH+46g6OBafr0M8aT5jUxV7YVgt3IaDSKjWhvtWhm56QBRdix/R91L29
RAC1hnoJ9cYc5Ikr1ip7KQ==
`pragma protect data_block
UoKxOQSkMLLe0iZHo6MzHpMuH8J/6GyHK3c7dUzbxDnV/TJZa46iARhNaq/Abyz8
/g999uwM0R2qMPo/GVKhWeZ1feWly0Q5EE6j3Jl8Cz0naaRGfPr9Ig6B/oYA6DWg
9QqfTLNWaFtvRv+wXU4CsVc+ydUKhUwMow1XyV6NAWsY1oeMYnlXjOaOPNIXQZ2x
4g+GEeBibpkHmhFrY2ico+orZWLeSh6b5GPP7ft+7ZiIM7WQYs4s3EGLEUcf6ew4
Q2kzdEyV5MDs21vQ7urOflhwbp2ZaVCFjBZjXKF59qjI4IfWeZJI3wc83nndbfMY
X6pXi9AlpnO37m0Rbz+Wgsl7f2BCZAJKLEFMM5qM1EP4lL/92A0eTDaAK5VtTMlr
aAbvWtB1xa1Rzjb8LIINbixvEcfgArHp6kpOt2XkyQMsv7eSvsUR/rlpVU/JMnO/
XSq1zD9x7jfKwre+i+872OXKfLuW895ZQ0SFfnb30Ehjb7nyPWAkx7EUgVQHKruL
9r21w+lKdM+TrQFRKZYl/rezDMJkUnvUkX5k/Pr27Bl7K8hVmn+p/A3ED3UVzm68
vrsRAE3TSK40CDFcEf5SZKwpkChq3p4oojoSnbfBK7SAmFf+PbwzlSWR2CmgjVYa
+VJ7c0gKfGsLGqsVIM/ldwJ8H9qOvEhINgWXYMCgDjqBXKeVzxaiMd+DKLFKQpA9
nELhWeRr4m6CEzWklwbS6aGfasrdQgSVRFb6GSJecc9tdzhOtHYJ1wKgw6qokSRV
SVzQgZF5YeLGS/vT0PNjNzpe83U33Ts07TrKz6EbyjqEBhf3UFLCRbnFyrC8zPw0
yA5OIBwyxLyeLBKo1X6hhV5BIbfNslVM7SWnZ7kso8dasp4qtbpXSsrhl8p9ePiX
Qbc4pjwxvlk3BV1c/vLQY9awgwNspjj/v8EYPWMkD+KbRV/woEYv5/xTeuHdXvC1
OlK3ZnsECuBMF6LWISR8MZINh3rzPz7fAZtwkncfvZUKh0NZwFShdHmoTTNtx6/l
nB41kvtRVxqmPzk0FvdyK0sFnOvOhQg6jt/LM24Nlxdfx2s03IOSz43+KhWZ1Pss
NrpMjEH7z6U8a7ZOOwt37AZMsvHuEcfokWq+R6ONwhiN7ldujtwoV79Rho33QZ0y
Ev017t+VXWS0RnvULWdOLA0wPZ+WFvfXxmL4h3N5/hJjJDt6SB2uuXhs0aSs/D67
51h+Jt0XtjQlp4BLTVESuNHJe6ATtDMLFwlOiJel26pep2SQgALLtwIP46LMq26w
OOpogx37GqsNWSyuX9B3X43WnR5vteMBKiWrQk8e+aWsxNrJwE7no2yVrOeAoeV9
I/siklCMfrae1TEV/K1qOd2MAo1aA+CCyAPsDrvT9DDKj/+yHZVHlzFnMbDs3xAA
0LWPVHKWJNyqnLoHbgFozpQTQzXw9sVR19RhRS4CYnCpXBSQ36CL1+sLbFWpE2wR
GhFe+b/VmT4o5BrPObyxMtE7jpEm83AmKT3ieTndKGU4gHmf6D2U0jwxTa4I26Ms
s6yzqa88bv+v3eGVuSPyYuDnPELlHbQeH6tvIKfIgCSuwP9qCBOdPv5QYQ0iA74M
z4NAdotmRqijLiVpXok1PG5hypmo9V8ABtRlNcvYzk1pFxgzU5bEn5c8lKxPBbPr
QrrVJ4S9zLkGufCZ4uSL+s7EDG8rAHvU5dskKQ/6/Hrwew1sHW7Z0TRZDNY2SUv+
NbmfyNMmJ2Zx2wDRbSTykn6o+JiVVloW8o6ymSfv+ZOIlrPwJVTwfd7Jo3kFjUUs
3/llqSzRaCsxXSdNBDoMv1ho7Yh2RJXmP5ysvQIPBkoj+XzjSe+admSoqRSDhMlx
x8GlAe0z/0jJ3kk8dZysBMD5Ye+i+8yGzIL6RBtuIdk+r7c3+FwUcikm8kRyfwH0
TIJ94MslxS1eGFxDc3qjj+Lu5HtGZakSVfGXllJT0K3vneovFN3Gbg25fF2bbtMc
JR9xQHNbYB2/h/iNreS7kfQ0S/mNPnW6QQEXd716o0diDAT7tdoZUWsD8XqsHINP
XIA3tv1m1lrdFk3Wb8cY2QrorRjrk2d+7unISpScei4ps1Z5tLj7rzLKZRlLMXrd
DbGHwlZVGF+pl+VKxVUSNtCHDd5AHOBV2mtAFAd1+b2E7yMWkfLKCaKnkb1O5NZZ
0JUHj6lOTaPo5ZWsdIXrdw6b1CLzItrX9AKwvR8Aii79Wi2Oehyx7B8g8dbJwRtn
ZzoJ6QCryevd0FkjQd5ktTVg70KStJMFFarHDzMRSrnd2s4tuQIGThO3N63IHTyY
XHooUeOxXPQpred1AyWtk+E7EJ3r1O3tPy5gaeQY0+slZQTwj4hcrO4xOkPXJiRS
ZZz2GsRjoAQrVoBPu/G//2h0YVRCJTzHYklg5qY4GiJyIqdycvR1G1ZWpG8OfVeK
HL1ZTMVeKfnfMHm39An0qJpoEI9HKoDTui85nxkCR6Ayl1h0yoH4eX/X3/i/KYJD
MFFdDd1FT5zrCkIhggF0lElccuqoqlxMzFkb2BQ/JrP+2BQOLEjKp+swCbbiwwxw
1Vbxj/Ctugy3hOrNucU8v4ZbPQmbbfYXwdpmuhAdMGymwIv2PqFWLOyrmy+nAb7y
9ifmtVbuaoxlZw2e9ZJ3CrDKh424SfkT0y4KwiXkKA6l0bQ515GkQ1FKvBoxfl3/
VlhbrnR627XXYThqFchWxPjcDzuzeF0LaA+bR5OwRoxDzKSqvyTRBeH/FeKoYtNG
R9pBnnJGQZR0jEde2MmpLuwCmUEV4+V/stnTUxJKAZzxjdcDxpq9LDSRnz9IO+TW
3rOyiITqAO779YdUGWF4g44TI6Uz7IAJCxoyrGev5IhP3+tGd/zyi/XGfSKDJISU
p7UaU22Sik6CsVvkXBTiz9RdqfJScEs5qOFbKMRpV6uqXgq+gqhub2dmDFILu7PG
3UipcMgzzfn6+5Ud9t0IofjdjlELFNvx19dAC8ZCOm8huKNOEvtk9Ujv3wgfLXBf
TOXO38sJaFsSXNIYSxNF0oO67MxUWDUjdthiMge6HGQ37eqpU3CF79fYrHP7ZPzb
hMFv9owTPx8Wkv0Z8jOaGFrpjnUViT8ZNQceJUL7S/nTwk4WpJhiNztyKv32GD/i
/88dpr6ZHuK/JYUpw3ZRrCxNN8Wu5S6NarC4d9dW+E7XzHtuGv+AuA0RaeHJxf9x
dy3ZUAMZfhh85yWCRXtPglD5+C5eXPA85pnq0+p2f8B+eKYrU+dC16pjcF9FekeE
LK+9ThOFRZwipaHCSvMOxb+beqnomw/H6ePFRJrhUDVrCc3QCTJpjKhEUGue1WXu
eS7inVcIPo7E9clxTJgdOVTutHve24qvQ8gpNw0H4qxg+QJ+dTHZlXWJGT8p7zMC
ieUoswmSCLouJSQe9YBB2DRuVY0HipgnDeW+Kfo0hZoKLQJPXL/IN1v9Rtp8qUUy
0SmT9vwcFSy/tvDEx8Liv7ONnBoWSRkHZX8krferjHWfoIi2pomSzqibAaEIE/li
PMM/hNzvIDreX6mOK85cjE8brDNvEWkix4RXtKszUPJrsQ+cxRf48TKNtm1SygIJ
fl7QMnFx/KYSFRBP/RLCYv4UH7b/0kXGFxrb2NDZFONC6prImFK9fSsI7Jvt70yg
YRwWc2UIR5ZiVjJKk6mI5nYukCU42usDRl92SRQK9gZ6Py7XvbhPoquxfxEJGeyx
TY+YOn5hkF2BqC35At7NWBbCr7vVptB3MSy2h6J8WdboETGF/W/qOpLsQi0d4Hqo
io4xZrPBpVz+cT7ay9FRhh9mhlQj1mCIe1/ak+zKQ4iZkTrOV3OMyJDb+2+lq8U0
F+EdxNNPFnfmVQoAPxH3jSzMiaF8xlWDbzuUkj2Kd8Lw6Uc+bV/FN6sLpnUFhMd2
ZMSXE0cHQbb+OZO4fG54t98wHEbG5TRDK103/oXW/62lh3vEqtN4rKHcztKkmJfK
1k5jHMeQRAZHXxwW2HvfF4Bf0RP10q3BVEscsYKBEFzsZ04Bd/GgyFkB38TRz4QJ
4fdbi0tDAUbbEa7lWbLo11fElhdcwMSX6tDmgdO7/NHx3KF+O/81Jt+lfbYk2gPe
2VuInOZSLrliNF0jbKVbxna0m+OL4hDoHU16Z79DQb/jVgQ3FB+wguf9kYbKWf+V
7NH+zzmeq24+PCwTMzL/Ef1sMpi8CgYm8ABylfa/P8M+WO4v37vnVlvkRED/PQ//
qKlfh6JxMDqOkYqfwJq7feb/Qm+LSLj2qOA89xj+/yvoiS/A0AxmeBjcw4BpMT5I
PUoC3oSUHsDbxfXL3zKwwyn0vW/1kZH74GIBvaIJVIA9aUVQSrDV+0f0SOEmaXbU
m3gR4Mq9dR3hfr9eDaHmJQ7tr47z0GcbtqubaDbXAKZ2R2huRA4eo1X0P7uNU3F6
9hv77QGqbLZz7eAdQXqE5h6utKohT+6lmhEmIMsJrhTYHC3RP2H8YtBwRjWDmgym
urEgKm0dAGMJTJojWlnGa3cnCjvOoY6+yda36k1RlOt/ul7P/WGmXcJ/LON/GmQh
8L4pAmZ5pZorINsCkt5BeCVeQaULz6uW9SXIrz1UbYJbxSYtEVBYtHs1f9ym3YpT
2Ak8NU1bZeb+WvbFdI17rsRfRLUB0pAdm5Qk0qJGI7qIDVdPAETA6xhF6ZhKL8Dn
NY7KsPR7k3D/Q8xCpUM2F2I8oY2f3X6Fg8oAxd7jqCnW6F60j4lqoajdSpnHBCnq
FbPdLfk2pXI3YNDbbve4m6ielqidrSGvEodKxJp2kmSvWzMb1NGa27ebYi9gI8Qp
ScUBWQWjyAVD/Yg1MWq6YazuvG8d5joANUXrEb8UMhOP+/jJYI69YBwYzItWy7l6
I7y3HoGcshR45QvfA4uNe9J0SVkRnUqsODuR2TM2VSep9dcLFAdoWp4ntCaBtElV
N/xJ0ZSy1lMr3ZWZYrl80OswYsvj/2NOYfjIxTUGGkygC0VE+zNkFaP9+gQcrTZN
gqQiDlklBlu3lpAbLuDOeYphR9+l7itVmB+PVpBcLe29bxmaMqqmkKyPC/SQ4Lt6
yFFliIQel+2AEtHHojUMQYSQMmIteleQAxfWia/YIOQ4RZy1kUhf0RFP+3KRqaKa
2bdz7qXVK4rdp0bqltjIZGBM9qgdWNAAvns951PYQo7kkkkwoERfFZ/8jvp6Kj2J
jbD+DxmcZSMy6R26RXjEdcU0ZxbC1xdFn0RopUk90hRBI4QY9/51StBfpnEIFCAU
n/6tNLcpOgkLWv51t/9yyhyK4ZWDzsrtc4jTIURjSN2s5ljS5QK8qcDoreujx5GO
3IDhPH4NkVj6ajgeENq97CF1YwSK4gI8JqhQ7PQFI8HRCPIKAolY0H/oRHDEyeIW
y4nEURBudgu8jHTkHYSGBsOFM3L33pb4DlPf0cMppvUhZ0hIfovnM0Er3llo9TEM
4nFUY6C4eGZx11flbguEFsxg+ADhc6zhVuME45TEhCDzzPnMqf1+nkHrllyq+E6s
dBkPJWt2CtsN0qPtZ/Jo+ijx0v0xrsiEUH1/PRdbopd1H4wYikTNwixDqwx9nYRL
FiS3/OhdBgV3vT9L/LDQ7Dwwdinl1VxXNilFfoPcvLIll0Py0BzjDJttKeNhxCjG
UCrBCFQcViTW9A2KgrnRIxPIl2jZxQjJHqxIOTzoR61zdMjJ0G9xO2s/wVIULmQD
q7I7S/GYjOHFNgW1nt6Zk2fDpNmYpntXs/+Iy27Uqk18EcDHrOV3nOXpU+USgZxJ
LxevRJ2FMlWCs1Wn27upA60oA64zFSYgPvZjXaTgtd3pcDRDrB/tS9tvW7p2IkJz
Y0at7V1OAQewJ+kdneeJ8sxc1w63skUv06ylqUj75k7P3Ppn86TtopAPLStrXIXm
y5F4ZiroWwjRbdvwgX0u80H+KAXePh8cwmYE7e8BZVmQrtC2JzEYXueNQEiCm0Kj
Xgljvb+XqYxI5PVOpZADlgDn97s2jiGtMBxKa73J28/igcBnHZdz8h3NhDzKUeTa
i7fL9xfefmGA5POCDuT6de/5MoRUWs9llXtMUimqkGpUAv9Jxd1AqiwZZ62Ru1M6
h0Tgngp3ZVRIAvrYjvitKDaak4bqZMc0YbW+RHpyYt8qTf+E//EJuOXypI7nKHlC
FzdEZg9kuUTT/qCbiVK975Ifho2YngzXZ58GLNd+FjfsFSgmCli1hCkGQDFG7XS2
pklD46SUMgaZc4B6m0ox0MsiTxMo56YffBtuxy20GWIuHldxhv91fk2Dg3jnyspb
2wBeTM3Lr5i8OYIIum+0BXyYh9DQ+Nz9moSvWI73iymAv+qbPgux0vO7jiO9TZky
MNb9kyA2Lkmd3JhG3tqpPdmhnpgGbcsdgD4g0Gy4qi1doBUe/RYrH7TNJUgrlRGF
sdXKcPN7TJ3zx7MzCn/Wc8/SUrr/M4nYggFi4xroF5/AKHrW4I5faq5Qt1IrQmQa
BW6gcbtPkR0mlFFIJKLwqgLVg+sU2r8BMEFGGTJ0LzYYP0VpafGD9ED0fSc8WEKU
IZMSIAvwepS0pC3KD0jYrJz3HpOkHQUQ08WoHKeZDz01RUXxm5p3znECXb7Nb4DI
6Wa0ZrkrGXsAsxeyo6JsbtDJkejws4tjHZnVBZQbHd58f4/aym0zvAkHGKthzFvS
N7hMnbyPRi9ITIcnxWR8/BBI/U9bavlaWp65/ja7egRRSurEDf/IutAxyexsxOm3
rbvQNEv+ZhObPydNNMV5JgE3pggLp9SNFOvjxw6rbD9b/1B4aIqDYtV/Cw4ane5n
LhrjN/aOHFp89HubZ7Ix+XSKk/wn99VEyPjyZfj2prIVbrvvakbf93SmyUAeDcaK
G2hDIJqSDwmdYSNldb5Bdz4Iiucpfxzdotb2mJ30U61o2MiYFjHpjDCO+ca4zCoi
eD/PSDi9NuCw1hjPCwSoQaBDf5Wna5MagxF/lo6PHIOcx/ruGOZgOyJ5Z6aAmK+V
xZLNTPU5MUxHAJIg8jR2W15QbPcXC7OiPX7uQ0lLraEXaJPBcv6oWj4eUrz2JvRs
WpZlVndDY1n2k25cQhRTaVzJUv9KIY7Ps+IKDcnaNgA3//ok8GhBnTLR7oB4Ud91
qWOPQfRTi3ZkMuYWQdIk7DgPNMtEapT7n0Xz/vxuszi3SWpAtdcLYDg8WxhazwPN
6BOVLLlvJVe7eDK57XHUpMnF+kic+S2ohiO5+gbyGCc8DI8tfgxALgnqjrRtEuMx
Rqe/hGAhSCTPhiYvdxkdC3jCk9Gfrgja7r5ueDd2HAonEzJRQaDYrsY8NvQJtQ64
lCLq6RqCyjG5qkLkT72b1n/PvIw1rZHafz7lLfOrl7Y7WO01RfWt/2MVdumf5dq5
Wl5S82aKPRj18YVuyjv3m6WH1D0zTLSc8jmA9Rs+OUEf9MAGsGzH+s2KWQ+E6X4J
55VF0iVKG6jLUyu4pvvl87ttc/5Mft2/DYQYQRMzjeSV+PXLSGJyXI4WKFPj3Rt/
Y+ZBjq7UOZuy0gSRaHNEK2g/FgYUhU5GVsGRbhp5uV/0h4WbccYbjIZThmfljxsG
cvJAIuTyaYXZ8TtK/i2OcL98jlUb5DuMyHSecaGI2pS3zZ9YKftH0wLfDrmA6CRs
msQwV2igabfv9pDErBdYiy4TasIetJoqLCThyNt3ZA5emEsHlOmHHIz9LkU8MrIN
KEsUevBW3txT4igyzfIdXGeoowaAKxJ9GSZ8AVxHzBDqFq3OvYDmGvJnMxEqsQAb
ioVdf6WmRwkOK89nAIPOAyb3HV3tU4cbe/EQL0OSCJPLzOwoM0cuJ5XKExcBmd29
l0XD1JXVYRwoSE7EPHnlgaHg8NCRUSmVxxz2Q0uWjgkqeJj+wAOkcphTaF3aBsAU
oW3fsoJIoYKl0Yok/Dss7KNVX32ilFBrbempd8eB5ioLSz2q0yXRaeVkHLa2EGLf
BZq9XaYAzqaCvgHlU5WzvfsPABiTpeD/lIcBzWDd4LCGVvklY0XnEs0dGCbrtX3W
/szJ/v8yhqWhBHb+tT9ewhyTomrp4YXhM71qmiSAt2LW56y3yDfFlwiZqGxNbS4K
9ANP+IJSUiK503nENgQxVOcvwd2wWTMrjmCUA4aatZFMWatBTn8GftouJohMRTpc
ClJ8ZMP2eCMEqa5vS+qhn6ETvIA7N2egFlk5tc9L+3QJqYrJgGAu9W0AESjtaEhd
OyApj6KOxBdN1prl5wN84MzmghiQOPr+L9OePzbOLKd4elpbXPjSroS87Z9Ecliy
GISqvN7dpEWLVAi6TEqTJuBwYfYY2IMaT7+TLl/pjyfQFXF92va+pP4Bjt4CIlTl
aiZyAxdFCek/ccPQWZqlCmu+OdJkYsaESAMF4GIMlvM4PJ+/UV12z7vbAQhxgjWY
u95IImu9uyJYjbRvmCgDmz/fW3xXKfWMzIBmB+SypP3y85bKlYQJNuYquN1ko074
cS737YgyMC0XXH9ab+7DCCXIiBqMaM2kr4hb0ZCAPu/45Xwloim5jkvDlfF33rUx
MRjpigGlTr/0ihCV97UOVQlibDL8q13ckPCrx0LdhBNjD+XhosMXke2z/dloieHj
SSwwvhUZysQ8+cr9566+po8NL+9QdDyAC9pik2mYAxcGQpsWjB876bdq2l6+f0js
Zenv1vphjDEOog/fEmuzdkRETrkSBnxy7LknkJGoRRir3zNZofMFEzdRJfUPBYzM
v2aIwZV7HuIhFNFsClYVZO2VLa+6hcb+/yaU6XbtYnpHrTb+XOrMLjlaNGtUkykU
UXnx9pSl5Z9UNSU/JbeARhxMwG7oVjugm+BCE9bu7NKDayEqPcC4QfaQ6YbnAFDp
UzIZqwyuAj0sqULknj/gM06OHZxI3Jm6XiNC2x6b58y46JJKc77MpZNN0DIy8WjG
L5imhhCwVFeMr+2K/skX/iNGN7tKyNeM1jD9Z9mTjrbOez0SGCt5HWcG0OZE7vug
rTGsoIsfQXmX8k0rH7LuhQ7VCr2wk10lB/hMEl5E3i2oebh8/SDFUMQklCTQl86n
esrt33i0w/0cTYggqOvSgDS4hqD56evUxwfUGaoMkOg9WdXhwBcHGtPIj654EsYe
cKtc3jEkdEqyPBcUbnlg9HT0Zvy137kTlEdnIr5MQtJFCYcdJ0NXfzvOBjJdIFkr
oLN1Kiat2qDBUiu+lj5a10vuYUZ5ACep6uWTY/M2VAX+9lX/3v3h+KhsUZ1j3rH2
Ag2vqzFz2ASgnD/XdYMbNra6zLdAEjEpGrO4yLcjkSDV8+dDkFMvWLmN1k+xOi4u
S/ylkJc0dLl8Ze2yKiV3P50HnTM4TNVXLzk+O0FbePT56z6qRb5AnGwnFJQ1DYTC
CB1L0gdNEwlKEYtn55sjwVtQaK9T2+jV5wchsVv2gtkuYdy/hjLbbipZlrbqVW7d
PDd8RfO7txrHEXl1qKghibjBoqI94Ml/4rfFC7CUggoeimND1C9KdUEzgYEiq/lg
CAv+Pd69+hd0kgoYNaFe49HWUQ/X8Mmv8qfJP4PaL+OpjToJLwFvWRkQqB1RSZOc
L1ADotylrPEUSF2r4i1IKX/gxh49+idcGZo8+0DkmeYc/Bz1f/CAv6ncSKNj5Tmf
FbuNAhctncsav8A05PgklUmlNW7jBMA7EamaeCrsbZ72TxvbdcWyCnx7B9BbhGj4
bt/Fx3nqR7ytD96H1dKZb0TSSdkI7qjYu/PiYoKcr/qDvlB6rad0iYuUPM6fwyIR
pGQxxMGTsCnzZg+4bmowbpPpEGfMSNQKdrCJZmE4N9txHFKquVmtv3iQ9W8nUFPQ
OQxXzBUv2iU1H51OrVs9Yo8TSg2w+G6HrGKSNFiomCewxqmPCed7G7cl4MYVTqTJ
qhSzXo1hAOBBBp2gg/MXvxulY3L9u72LZtyciWS17JxoYTF/BMj2CMaKVtPaqqfo
2hv+TlkKHFuXflB+/YlycwcJ3IsaMH3c85fPs8yhL/mUzJR7KFb6Kwezh5ltfyGc
Xq51fLABIy4XG/GAQX+hmc+O8oO6ZupDsQRk2MksA4wQzfRnGMeQjZ+YMYSP6wiL
GIKnwH7Z5ZmOErZ3SqCahEceY3je2FNQFjw2LFjBsG8r+NkwI23X1PSktaKybewk
GMMMyn8astaVaK0dCwWKRXTip3botcbB8zdosiPreeNT3CGuk8I04sm5NqSX5ltJ
ltyUUbuocemLjbksChM4ckot2RT4pZqBEBoyJjC/pKQPa3wDt//KFIWkGpCVX3qo
Rw8Pz1WgNBaSi3PSCTdhQgk114AjsrLCwU7cs1l6YFSbcczcV7EGBcq2bc13OlTv
uDdAnsr0Acboy2wx2pANCraG5LWBjXO9eFlUlDexMIRu10PeeTLmJJJe+o0l9XNs
8/BvbtsDWRxy91NjjHHko/fybTu5iHlN6It7BkJ5Z/VH139E0Syts5+uRqAJLMxQ
bOz7430vcPQuGjPtEINGE3qymS5sZMvf+gCXJYYfk/S/k4k1gL/My7YIIROKGqQg
JaazWIpwG6IRHkcqBMUZlAuW/fdMMB70kcpz7A5sa7CojUD36oDIMHkBxsZj4xoW
B4FzB5j+gMlNOcVXeyfREkoFgEMxp3ieRe4dHK29V3vmz88C6YMLqCLESCjGcOMk
iZUNFocJyN7oLxH2xAUKz4FXHOjPLtFUQsYi5n48eD48ibjViEA+9puxJR69+odd
85Anvm2/PGHJfI0lf4h0gzYWe995JyWv+BceE7n81nKWtjV9GuDapd0EknbLaKv7
7qsLorsA5wQJ2E6D5HWcCZzVs6BH7QT4dmOI/p9Y3ollg7wErN9CMcAd4Wda9G34
JEr87cVnGAj7KHyFhFiTf8jSY48zWWGNpepgVFhLzq3NL+brUdzsH1EZUG58PM91
qYueYXRcsRydgpcDFanV5QwA8P09tcb9dpft57ahTesR0S5LLxvB+tY57JhNX6vE
MMDSN1PD8FqqilXTgWm1Tm5BqazWQAnm7zAGhOc2HiMa57JbpPwawZpBn4T+Ycxk
b8w11gMHw+QQYQYpK1sKsb5AlNXG9zFvGmG46yRzppCtCxJcT6RmjQWocMGAW8oC
9/9rJD9/+FFws4t+E+c3o90+RgiNW+1H5C8ZMDzl/qpdTXGbKful/kcJeLD+N3Zy
3TrJC1Wo9NYQ5XRJvXjOLR7xS1Yg2J90Q56algn8ablje0fqBSBkHbQHqBdYXZNO
lmXn2XYs9N2j+cx/DSDKhIOisoi6yY6labewLQGcc0eKkLg6HBUGtxP9oMXJopy+
SCjggb2xYr/9qbT3XzEGENHfO+nvtZygRuV9ueYwZPxpysxIAPtywyTe3AuYujer
+a4U7hNjMEEY/NIcfD9MQ9CJE1esh6/R7vltc09wYS1MHGGC1BEwevmfhLU3a+IZ
YBrInDKL+HBwL9ehBtNLhidcWlUqKdgBjIRkSen2fpiUkhkAvePrujTj+4J6j3bJ
R0B4GjOmkFAStLvSy9y6ZQd3VLxqDe2jIDoOOvERBkcSCz/nkdHICJMRi9HcwjJC
1PI+l2jAlYm8AUJvrQ6dDDkyalmMMfipHsRqRZJHbOYATTUfr3FVjX2QFso3YsG3
dTXGHCGhYM/FfHjRo8faPTFGD1ESJaQH6xXKbrB6g23qgz3bVPpqqXhAWlw+Qx5w
tTGXS5HUUjYVUnEhJE0B0/MaWZgNRlKUNEQn3msVI7kOv45URp/W+7symiEIZYVt
hDdU9+wyB/m/ab9Fc2bqE2UrU8Qjd3WFKEL/s+wN5Xex+KonUYIvgY0ySEhAl3zV
50GFh1pI5z3U5PQ9DEK6gFdUoVi2syByOMgwHJ8UAl/oQZjxyCW8dmJQLLd0jnIF
PmTJgLU6QbkX7GAWHld2WTNviC97lTQV9lPHW2/M5S7ekQnbmJKXlUgPNGwILGlL
ZcAGK6feKfeLimA777RTO1Rr0Egib6cStTd4BXeEAZmCXb/MHdxJDdsM1GLKz67w
0orQIXEj+mNUvZYe0kTznq/EDDv5zraWX7zSPHJf5Tkzgbm6p8wfo3EAdeUnY0Yl
FKzcUmPpY0g5gSFrfDZymCq3W1JVCCYIrYIzTeWzyV2Tnu+BWWE3cMyW8SdC4jP1
tMup4V0BlPacPiO5fVOKcW/ZaRtBoIA3lkaPyfgnEJhPjV3QTJ86XfsYYrzf4qgq
uRICrEsLaPT0GGA/UYbOA6/5lQb00TQR/IMYJ00XK/evSPcLABZ987FRZu2dpqLh
U3oEd/euLldco6p3msEj2ej7ciVku6odcjWHcG7EPSRXRYQzCD+NZrEvoDZlpvcS
VDrQGnEhdF/hLWwPFm2sYF0XMGzGmSfRN7qcIZn7pQ9nl2dD1WNE67Rwcie48FQo
k+8HvKuquaKoxFYVwFE0UlyAxvpjrKto7JA3p5Zaf+bNfxCohCLkZrZoeB+0KAU9
ouaoNSoHi7kaBccZSxnhbrYIvydjI44jalTE0ts7ffN7x3N4/Ay44r8YJlVgVqiH
tYHf1SKKXOM8xO/o4mJhX5t7is9zMTK2SYZUc1XQIRadOExV1oMiXEkgXM9wLTug
sdkIR3DSEfsLL9KakamXmdUWLtUMW5nNKr9ELMF5zMwK36lzeA8TnYbGdDsV094e
15CYsox67jtc4tKwIRqpipwJmnVYGPNGhQBKvCq+zayk52ycbYjSz7JgYHTBTkYf
Cc8altFDUYhJI2x1yKkdnBXx0bVo14x3dxbNH9WfU7hyinHFRshi6AX9aJSeWQZR
WXpyqwmon6Bqh8/5DHV4EQL+r35pEtd6InXPCqJtMZffv3sYjz2lH+k3JuGjWT/b
ISZbMAppgHzwrXm+Us586N4gWoPiEWmE/P+7Plx+rEPPz6DOFIedsJ388wOQQZ2W
dZNmgm7qEvC6F4bFCFdh9aqoclphUMemFCwn7MMYG35maIL/BeUCWK2VoVyEsFc9
aLwqGtP60uAKP00QsRphdG+tezhUrHwz9jiRCKxVqOiQA7LrvcjQSLdCLujV/29M
xvUMzc+xvUjB6JSyDwRgRS7zGEkPGSbiuPGXm90xZ0Dmxetrgg18XCu4Omuwac0R
ZK7ZL+c7g5npnctC4vRAM8bBwxdv1FbvXE2VM7bDn9Qzie0adNSr0nysyz8dLMvU
aIZwriVPCGb46fyb1cGQ/Urm30zSpQoeb1Yu9y8moOEmdbtlw4chSTRDCziABTa2
CXI/9Hk6gMjr0YSwvcZl4GfN1cb13UBKweLgT5aNMirNprDhjt82riPX3ebLL8ee
vxQApjCndT6cs/1Dh5+bHPayOTXYCbx18RBCeebEPdPO2YQP5LxFiXycqHA/04/3
K9D1vNmL9S3NVe7d7RoDvrI0ZnnRbPLlOEviPlT6dnSdmXLbVsOekgIqNjiIM3o3
AbslZBW0pK2HH4JkK8CUNBG6ZyEJHEJ0OeQDH37dgMhfQWqOB6aqogeFEJ1jUYWM
p+6ljSS5zC40vRx+Kpi+D8C4PvEcKCgdmU0kAy59VOgmhUh176AGvAGiq2KCca3+
H2SsQ/IozRour6VXQY3Awm6pKjxuVETy2hiGW77BNkxVw84/YIyt+ivCB0umJCqJ
t6kd3niOZ13vPwHTFeI2uRVSeE+f+cHeLB8lJiTTEILNniWSvUkOOgpk5ukpWNlv
L5EQ5C/63GrcNBW105lEmFjaE1HrFtGcUip1Rz2wWgtGctiPEn9iLGTzaDucNXSy
L/m3546v9QZuqpWrPv0Ekd0dhB1Gw7QkDjmLUkY2neNDm8pgobWDaVqyarkh2M9d
4WZ5zKiiTPmf74o8AyBzu5XAmOlB5b3+E6l/UckC7C7FVUXpkHdNSF9jmsVCvGqP
BWc/D8gwaGSK7MpC8NS4GCH6+pyfyGKUwc/bK0zQ6V2msTVUPXxh844GFqhkMFTw
USPmpLsa7OlrZetliKu8DUrhZAddVm9jpYS7nCkXzPWKKNDnbZQKBuCpwNT+ZUrP
/G36lQw98ATWgvmxQZlgX5QaCwo/V1rI+wmmF5QC1XfGGm9tBPowxXLpZHKp2k42
VwYzX+e8pOUGnRzLR+NyCD8LGKBM5TG7QuZct2xddFHRcgtztw2N+O6Ws+yX8B9h
2UFD7EneTjSoDB59AYfcIlzT+9Pxgjn1Pz5eeySzaqVMgxMrXrih3HpWTNR7eBIg
JRHa/t06tUyfKVa+WZ/KTkLwZnMgl4qLPOywbVpePmgtrfrT+vWoFNnWRnFA6KHq
NqfNjmLQnu+XnoQsWdj7uqQq3UjFqKSH7YFHGIjbU0+8wWZf1bRzwEwCT7/OhgSZ
CRKb9iE8tP3BYbNlk8FoEA==
`pragma protect end_protected

`endif // `ifndef _VSL_ADDR_RANGE_SV_


