//----------------------------------------------------------------------
/**
 * @file vf_axi_env.sv
 * @brief Defines VF AXI environment class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_ENV_SV_
`define _VF_AXI_ENV_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
NM9o/moOS35QqOlqrAPAQvBl82AMwoEWdSJOzugi4Nejc6ta36LfI5cmj7//B1ha
GvL94PLgMKePxwHS+/JsgMHXG9r1EcJGPkj7DwnJHxcWG9B5DdKAJCCvXb02kS7v
OemXAPc09OvattB+Aav8JHR9td7kUxiJQGb9H10k/h8A1PXnMYPaZtvF6UospwVZ
3Nnfk6fBgfqzwmi3zjRRtNEFCLI7BNgeH4HSm30LFNFGrmaQQvmvllzPzuhTA2MJ
9MinqJV4aFOqUeu2js7KC3HfqQabIJFI8RzJ2Q9exXOHruD9dTszBFobIMP4+5EW
O466ZTSezey9ivd1z2Bkzw==
`pragma protect data_block
YUFQmS56xEQXAciPPvhMoxNbMao+fd6Iuqv1aMXhJ+vjfAEEX8YAmcADxaZaxmI6
L+Lp4wYUCxM4ejllpoBLJE1bjegD9TRqifK5e2bGdDrulyPm5IZlzpUYWgawkNgT
Vtec6DZIE4Xe6Iw7kqjjJz1aJ8Z44Meqm2em8f/gRQUaWllBW1MNrrvqo0s6wNad
Y1EFajmdn31ah8g9fr6EjMCd4vxaQj554PHMertMJsXaQuo+N2ZEVppSr+iGN/6F
idKUNVNBrCW751tmy41vk9zVSa3PEhEtWDkhPdU0DICrbX6eL649slDHv2U7vaIZ
M2UL7MBOJ0oIXNJ7Upvi1ZSZ0fk/8kuovJemr96ScZ+5Yhb6g4iNUrMid/fFnTqC
vWAS5ABYov2lchpprNg83P6kjhMzo/iIlSuob6wHofadz2laBg673pbozqHnCXo0
Y0jbSzgB2d7rgA0GhJjGkVnlWdXX9RTqEKqO5uF6dbd+7wM7qYBc+RCooTXb9VvO
iA3lm2e6bwz0dn/ssTJQfIlN0+SWk3eCKOH/NNHcVNq8MFbvhoCW5JKz5YnRFmfV
yrSTbS5E068pIAAAw5Mj/ZzSLyhpLZC8UEIk7O/d5owZnZ5IrQyufZdxIgSzrQNA
LdFRBo4I4MB4gaOT5f6Is0mO0YOoM6/F0W/2NrK8mMtEQmaq+ylhAwH6NBlqVIZx
NSOX0xs078atDjhzg6X1KKUf+5f58ZRAMGdxCHCldYkLJDPKzZgdkeo33mRfRGjc
opAxr8DNZsqv9fvQDdrAMk8KsPx48BlWKQJHVT34oYVEVzHmoRmvLzspxzVgz89R
pvQrA4HrUdDcuAKwdnPxUKkR2/xC3DIJpjR1gQ1Dcdvfs6pdnq/O8DBfICwwznNp
4KMtVM0Nn7eYbU+3+NnarQw/mz/xrO3/hyrozKXrRoi3K/ZKYXiX/+9fAg4FmpCH
A5HJ8BQdKc3YiXfHJeGaviodxOfWlSn2QZc4/iBhVOQPfbeSGUjHc2JClKW+Hty3
MA08Bq0vLLDgVbmKKTf1lWgDsTMEsNIdAjczgV3YWg1goelJrwdbfEmMDKNJQE8z
bB4Wf8LIG6f+7DfuYF8m2DVPw5vki+7Hk6CQ0A0k2TsbQHCFYtV86gDZUP24BA4E
0dnROm9g1G2w0+4oClVMbTot4pg9hS/9nCuWZw1aFZKp52pVWc86hBJ4GRV8nwXc
fMdy8Ah2ObQ1347qBKW66o2l4mK6fJ/x8obr1KvkKXySO/y+msnVG27oX9/ztMus
rsMks1GRsixTIG1RQJIpJwDLbYJG3HcqY7tdQyvgOgxMUmx4vtoyGrnAn8j+AH9I
kczwDmennRFzoEqVeSF1dcUDH5QdUQSIoYgnLRAuEfSNCJ4sw++Uf8Kvjmb2Gq37
IZ7T8jxhd1HNcs8aRK0ihU3flRPJNifOU/JkDM4erDyh1hQlPk3aHxfBulIqH4UX
vDtSww6oSznu/oNJvB3k5YLZwWrbeMKgmYhyYkCWJcRmuoQpN/Z70rmQRYeJY48h
CVYoHSrldAylEuGG9OV05lItk5LXdwt1+8iHtRf102sFG4xGYnGzRaoDLD7HASN/
WOJP8mLSa1cgKZDvPI9e1x1IWyjFFSiRMitWLQScPP04/gozkT1Pm8lTrUFGeoXg
6uNyDKqbhlN3h0vhgOB+J9SN4r/oPbDJn8cav6PLkRtTzpeu7n+fGzM4mzVi34J4
2taL8N6+uwDxD7I+P4pWaxqbunn1QJhHk3DZoILUF7tWUjbIUP/EOJ+FP9yxAqx7
Xl66QZuA7onvjbVmWr9zoiwBJaT54SZoGx/gWm1jUEumpmVWxJ2e1sYmNtswpShk
6K2a2x1zsdJY/KNCYq3m11Kw44QQwN/QZKcstuK5xpKDMwrU+JYgNs5jpByEnDZJ
Zr6n2T7+fBmks3sI5iB8KjQeEblLWPEjZ4PvRzzuq04KmYLE3EPUJ7nZ+h9tv+lr
rSuSHzG9wrnv326BQJiOB/GKLTDZ0p2FAopHM6MYH12+tccj332s1a63tbQCdERX
rLU5Fzg4GRurXtljjFQD1QowuSEEGm50Ag8m6AC0SWyA9S6L6TzS8rZjhh5JccSC
5SoBIwXqvDXXgofB9se/NGJ011M5Usu/7Qj3Vu/jvWazpbbF3I0MNLmcY+hoFgLM
usHVXNnhgyjUbLd28qM2wyRCt/O/OXq1afqeD5KGIUwQZh4hm+PrFr4GL2YFHjhl
Y4YM37BhZZ/Qf85e533tJQvvvnrbBFWVCaGZlfW1n3fSP4+NYDhm9bfqhvSp0L8D
mlFIXxl2q1DmF7CLILjlB7kqn978Qg6cLbDzI6daob1sVIQK7bdzKBwROOXJmXwY
d+0K+TFKDQ/NFVCb7nGr959HE6sVXylctUI35jnvh6bDz4fzg3F37Wlrdz6C26DR
DLsIVxNR+HIxIxmw4nf/LkTHbUozOuzT5IQgR7NTulN3HjBITxKgoVwaeXoGrnh/
yUGc3HjzP0oFymUvznxeLBri0RQF0C6otyJPkdytja3drvPKQUkV9AOK16BENUxu
M1UzwF1ZjLzN4VGfCCdHgthEGDu+F/1XDTngArII5KPxbEfyrCh5YXC3AglgYRf2
uNdhxaOLNNR3EwIOS2CUhhvAI09rj35/YQ8Xa8Gb/DIN51BoO+N94+CiR7xp2+Q8
q+muKlxI9fQHlm4x+f90Svs3HKe0CLhkcwMVYuGVRZ2PWqaUGH6BZKUvwG7QE6dz
+85tJ6nLeo/GmEvFT+QBq6RF15Lo4jPZA6Crav4O5bTmV+4EU5iha3YHTVWVAg6Q
PICSEHTxsqAzfKTod7X5O9Ok9pMPljjPC1AlWg7Z3C9Bc+Z88qYYmLQVIPE2pSQO
M3axElsGqQ8fbAOG1GwpuxJDSb2eD9RJwMq/KK2kSydhRxW/ckYuT2EN2d7u6KEC
mR+EBANZQdCmkMA0f9oLIA5jJIKG5arGy7CaWJx5diwrxMXDrJ9Z10oaZbKUfcy/
5FPg2Fuj+bcbtrIRpyS8dGG7qNzTmhMugV9jbHu4yQytbvMmxbm7mGezvGgVjnS7
4aabomBVAJnLmvEEuHMzcE3RtluK31DQUAuWqI+JDuRmS0fOKqKZW+daAOYDYUBu
takuZQ4Vj1Dyd6zJ0nrhJunGh6Ao5H94Fd4fiQLOnoyjHdAApV6EBDzMhgE8v+P0
FQ7+5aPqBzytlfdCqGgIH3JUUJgz+Lqx/uhPAzebDImo+1yZnwYtuLMG7qoPmMY7
Kh6NikZUUKiUEnkXegNMj/NkDlRsq/kKIjuDsL5jR4mgsYvZx+TkRPuPnJ2Nus73
hqyVIXB/vrrjPzxOD3RmZin9QRWQmLpDVfUGwR3n91M3O74m6omgoH2AsyJp8fsF
KXzLWIoXqvw+kruSOpcgXZLkmy6K6FjWWvHxylRX1jnegzWROhgCQ44eG30qAgGM
E7thoG0BVeuLgl2189mrMP632gm0oTaIJPYaj1HTu8GL80SNEZZCPdPDgiUNTsHl
BfRYyTPJhZ/w0qRfg9vr5hAtqG31ICifWZnU/34XExaQonXbjVOWsGkY+rxdcP81
BTXkyJJdoZtD/pqzByvMa4uAHTcAMjGgOhxBqivoBNo63goweM7jtL0LSIYIfoGL
LiuIbp7f/+TSyGPeQzqF/Jik/bzXCj9DiMdUey9UHcf5KSW/zaEWY/EKaFmvggsA
SsyXaPeElAETqngpNc0vHTrS/Y+07mqxBiVdsQw7QKH2+hL+8ydLip8TJ6++gGIS
zNRYiy7VVQXAUu/gMRJ7GHqww/DHEEAZyAL6WICpIfW/h2FAKnBxra7JFa5luXZn
T3hKMOhK5xv1BR0dK+y0MuaiFvPiDHFHRFvqbKb/oJcfNAQAjKWr0UPUNVDqzco/
OeFei+CRGfX4R2JkfR05niIqFHag7CLW8ckcCPfpEJdSoi2nA1sA3lxsXZTRdyM+
FLzuCBPVgCHq0QqpT5B4oJNCEcUxpwocTPy0uAZ9jzNvQcY9AOQjD6sOxLCFRw6e
3u83JauWrhxFfh7wNeN/1NoJB9TYMGx+w3pRVs0Gw5O8ofOraZ70sA2qQkRdVEX5
N027HBb7XSbAX8JEbWDs8mENfIPyANC2Jdx6M8c8aFBlsFNXo6n8TRiiw9A9wLoN
NzBQLVcU3sabmz+aP7xTvm8csRJRg1zflPunIHSM66A8KfcQ7IH8TvYHqNGktons
sorXVj9NnMi6tzcs/Zx05zC8QcNEPxprKULiZfIPIfMWSEJP7jxmbiSa1fT9YHjq
GWZLEciPuIUF+GsHOqLkit92ZDcWvl8bNuNak63IMu35GWHfp1Jm5BZTT60JLXTQ
RMnGKSNaBMONkbmn6oc5RY1i5u4Vnt5obl7R7A3IBQBb0ozfu5nGDPjjuWbODzKj
YrRp3sT9xgO9fHge8Yyg4JlaZZIhhzkMOh2t9vD7ngnTFdfWsDL6ohrkN85luYz4
XUTDfSm3PAQ9elSK/CCc837nyk3F0u8QW8e1SRsVy2RURuYW8Wc+p2GvgTc/yEf9
hvfCfGHZvK5GmHY4CtiyGvRbozXSplGtWsiX7vEydH+ViRr0BJSV4RXe2qDDEdcG
OJhcCv1/w7iW8R7+hd8QpdI2/ntWZRQmKeKP5gWP1GoYqPaqc593kSJ6JDf4SI8I
AbBpC/wcp8UJxUVQvB3khheDHjct/3sZmhUgmKbolEyvc9Dok2zBtxKIBFcdZmOh
G1RbqKi0aVbpMkR+Q8cuQJjoP0JO9/ZS3HtMiOF5wN98O98NilN7TQ6cBH7tqcMF
gJ36+uX6hNFQAsdW3Es+mCd6Igpqn+ru3dRkoTk07YNf1bSdT5vdKS66UQuDyQS8
yvOPxmgN3Px/uBODA6hjl6ItBmNhrTUUWm6Q4spZvt3RLYzYThebB6qP9Hd5eLkH
upst0ClAI5OcUXvZO6cUVBKBOaB2TjrkH289emhpOpgj+7P3LtT03nGlJCs0WP1x
xH9prOI2guTKWDc7hz912DrXaj0kmrRiX/j4RxXyPUyKz/uEPhft7xZHnY31jLjU
mYqjCqlHE3fSwjf5D5DOfqoJgaLzfKqGdPnu0YmnA/4vOmQrRYPQggnLpuLNbY0v
fR7lnyvHryGFCHGjMBjqs8hcy7l5gdKlCj4v5l43Ohp7lKSckef8GAPz7i8gGDdb
UWjONDE4ChIOpe1aErtQk87bQn3kkC5uuyOWERv5VF0SzMfnYL9tntx2ZQzfgoVX
G5MF+tpiXWTzm0zs7pIiByZX0zJ69OiahzjB1XAzzQPhhzOMq7xgtwJsFLHIp/wv
OSK4R5Rcfz1ahLFRZylSqayx1i3H/+LrjILcFZ/tcegi9Pb/b5iOvHIgOC6lr6XQ
JmjS7a4ePp/kFgbI+5FWlA/wVcmlQg2VaYamZIXXiuAYzhFwhXbon9iAFMyucrqL
MHn667IW7Hw6l2PoRdbLfUxl414AU+6tqZhaqsoOMtvnbGNlu61t4F8kydPCfuBE
YngUy0kxcew5obgrj3y8m/fzxyri+XAhm65QVWhEpeaW9Z/nL6XctMSU5q6lEurV
1L2pgYQkpg5zd8BmNU7sUrL3YWDcO+9Rl2xv+mFiL/kmm77IRAf2oEsknH0nLkGJ
luieJ0IvBEYl9Rqc0LuD1fi4S8YIxAq6pDIGbCZI8myTEqqbs56VyZl2Ebvby2XH
Buw8nUW/LeNqot//sxetHAXzwLtIdD6tVFGjOSegKgIfeprVFEWHvYGOcIQsIZch
8cXk1XVIVAxm9P0OwG55fdw7BjaA0TETTz5JO7dtxKa78AMyG5hXu+5S2CASf39B
lf9xOSwv7NyZYlfbxsBfkLanX8UyJfQX3WlSFjK3TdxL/hf9U/l6K4ty+X/JwcSL
S0oHC316ucc+2a+7wV8jT+B2Xv4+B/kZdr+XP7dBhLQzk9F6L0zEmhndGOi11JTX
gm6BFHLpEwXJS+mpSluQMtQfXz4dZq+UQosLB8QbY+tVKzUCHNmxJMFNBM2Sr0v3
L2t+qVJxLf2rzx5ndiG7FzV76yoIKr1N4zUCXXL1NY6JlXLA4Nye4uum/uM8VhgU
ijgKlCvxXhB1V9TGEd2Cxv50PSidoFGVxh58vCBB4ZVvYWs9JPUKUxVl7iGnLvM9
5X3Sy2P2CrQht5sN9xn0dUD2xRvG2Svj2bT4X0I99JV8AIbyO+VV5VOa3VerHXHz
6WEqDu00TN4U5UcoGe0M23KPU6hzM6zzDbPpgvrRi7EvDsipaqkd0gp3GOyveZNP
Do4dcZslQUckUnLQ2nJzaGrqbLbeAZrm1DulB+0XP9XAPWjzr5ndnUCn7ZCCSMRH
w9HI6E0uUVJs7iBcBczrIi7d3IOx2GjKiCq+rLFGyQ6rQYKVlRJCIP/NZ2oYycXq
oWscy1aztptGLqQ6A5KdKNbgy+W+8mUGvGRaE3AbVZpacb9ST702B/l89o42inMX
9wMPPSMLWwj3X925sfFVU8SShJbAslqMhrjBvhgZAoK0BAE2WB9vRG10iVbrsXpH
aqgG/65BG8YoNaztdg0z3voVajCrQTunIbA4qSr52vClGPNxQq25NfLCvx+l6BrI
L/hmmgWi8nGkIulhAD1KL0KJKLIYXdZUP+5PKgZyJdzG6HdB3uCElH/aRJs+Al1X
B+cosIcI8VPuTFqkOvaTP8idfCTSHBQfmVuCfcDNvnLB2aEjlwzK01Oh8vkYfSNp
AYAqUpISjAQv7vGFZD2+/WiZvMmfBbyU78kkwe5mrkT+Kx7DRefMo3u8plTmBY0U
ew9hBuCGZx7Ax6DC3GBaT/EGggvRtcv7/qetx0IFE7jHMxNGaxK4Xms24yv+o8fb
haQEq5ALY9jsN3WrHeWnmgm+8Yuo9v0qwFM+cY4QSdjgBysQPm+WkWR9Ka0N0+rN
5WD+oJBd+NKejAdpMbZMSXgUTxEptBJw7v5OBq+w7DP1onEkwo6Yz+xO81bVxi9s
TDxdYHsiFxSBK+CgYslfa02iA+n32Tlfjg33g/cv17uOLS3IVCz7aEO/WxPV+FlA
RfMbokxAm5ekV58xO7XGtsgMeZuuNc91PyZaFJa4w/6zu5zTUdIUH3MLmMcskuSh
gZ77oNaAqJUBnp5JqmL/NdOUpWUk7dLZuSA6ojV5rk8lHKqgMaLNwfhFaVUp59qn
RPUIiTC6hjES+r/RCBvsOT/zCIfeAL3ojf8hKn2kYVtt0VBvfefgPm8dnH+NMkas
0QP0HExM/3HqGsN1zNp3X/r1ApIE/7PVoHCqyR8ZHgLE20JIOWYdND8br8eiznn/
qcPN+cKNtoUilTRuUDxLvv6g7/FoPTcBmWW0EQmrTHqRAtf4xnFd6w0qmdxavfOQ
LuSy+Hc/XjBSstzu4gCry1os35HEXTtqqMZTX1v9mrZdlJGjlyR1PT4dY7EI2+RM
Xkq9yte//SmIYocq6ANbXQcmA0vZXHTfYUieXhqoE9yysfJKbg2wOClomFRPhWCd
9Xqu669rZHYZf4/n5AghnaT86EK2YzUa2OuYMN22kI8LagkJFebPyTIVN28prcfT
/ZGD1ru3P3xMq6t8FzMMh87/5V9a46D13ImtTdxczsnFOy8p0fG3zlgT4ienPbbp
HJzjHoW6c/rH+ZHhth+i1rWmsMNGJarsAx3RejLR5vWPWuM0YUD1jSlW3sML1Gdo
W/Y+2qjUlnlNZK06woYT9m2XcV4xjW30388N169kmRd8Jd6Z9lw5B/40QlKe7xau
BXkI8RpJ1zdTIfJ4kFgLNmH1vVFj1+SrmdpGtja0wemuW8WGPjZZxKzPww15B5N5
IM3+/UfIDN7SeTH2x0wT9nHZP0LvyHwitKMHHV6digyCdbYo79z0GrBGhYiAXQwG
SCEck3pqb8+EXMo+0RQ7M/cww3uvaTLuTl+iKKtK3p4NAiKOyzRkltGQ8mNuNMbD
H+cHWJuEGM6dubS7HXh2ZHH+MvSS+vUOhITZ8TQ8gH2fQWBdT0nZwjK1ioJGpb0Z
V1bKbN8gBAJLhmXuJ6J6AusiN7tjK0kgyzDlHCbdn8mV3xaVKREq1V6DIRbu6v6C
odyefurmN3FIC7fswn/ObAB1bOw1S1zg3r0Yti0JLS3PMHvfCJdl4/QJSwyQL4n4
3qYv7iTufipfOjXzWKhAIQPwPKvcnkfoA9k8q5DFiOlyZwZ63ve45n9j86ZP0Oq2
fBRf4Eg2YpKwQ3Xkm7hGGEq96wOjMH11GMnpnh0Bmsoa3ksAfxU2HeO+H+uj3p5f
qP5Tov+M7+C3rpVQMR2JJE+LerVh+1p9KYzs1uuMKY9B95m3dV92vMsRsVJepvLO
r2d40gDJv3otliXbpN/4P0axvAGrwxhB3umflVssIuI07GXyAQhaCtDpHdcXCMEI
/Nk9nYc5QlBZ/1WjCaOyvJWRdr/puAbCv7/Z62jxZV35DqMjzDL183WT1kF0JR36
A6SKcneaf0NzRDGHxKFMve6RxetlGh5gsupDgTuwgpbb1KqKkRCsYWS19sLkWfeK
y+4IN41zQs1QBo6/JLWiKYPbFfqKWsXqMFN9ynqMazIFLIFcSgXG3F9nJP7PjPq9
sWlHjq2YuQCWxWR7scBbn61hqonDbuqgGIFBTeyeZB0jxTfOtz6v/npq+Ta9oGjc
0/yUuNFJc4FRmbTWRGSlxwc/Gu9jdlIZdW0He4Xgl9qQCLKHrqyA0/3ZgphbKs4g
MMS+CTsFYvskNYuCp8an0HT7Rd8I5Qa2AnRE2WPNQJ13bIrlBQoWWlx8Jgsom/v9
xQe/IkM6G8bkplgftPzE+KPYgxXLsRIFiQ2moaS7GWKw8lCbitxQhS4lfnRa0KD3
cnNpfe2k/VvIOLeMAh9B+Id/QBlHr9bJ2bEcknww27NmDWZfyJrUxjetdkQLACpA
RLGrRi5G0Ixa716heZ0oRMM2epSk0wUi3YJyhTKkMZJ4Rjct2RRt9NoN11o4EQh4
f+T2u9VqBI2oj2SZtia91lXpM5J9A++Vn6TW+/kugxdVGUfwROfyiiMRjuLniav4
jrcdbrHCcR2Wk1jdhJamVrfec0PG4EVI+O7HoJKhadDr+9WytPVPwiT4diyvz1dR
WdpQZU60YrEtESjsDNemDzix5ysWx+zViDbR8QBENxcDF9MtVNA6+utpdS5s+JU2
lVERoERJ2s6QGolt36X0DW7+ErUusKFoTqRMRrA8+ymvUKnWAFhtQ8wn6lJZCBtH
A4nuskrGTR5v25mBbJhIoYj0n/eHhmykJU1vmio51oZZ0IVou/ZcXUetIewMztZn
WgQbYloSec90cPTM0NQniHerxPDmstInkoaewH7UPjKDTA6Jb14net6vjY54soUZ
+yZOxeLSx6I8fV+CxTbLy6U6aciK5hQajhsJghWpqnDWAxsYw3VlrA3Tm9+fetlV
vyj/IYBO4ilhD7xmqjDqM0RznWtYgUSgR7bvluV1TkPOVHWmb3FhnRWZQ06INZRy
bfwLdAH5lB61RX72DkS506MPiHLwj9jbNqbZZWwwu5r4ZsojouE2ZSUSyrY5dIeH
GTpf9cQhQVPPLmZUxCdy1Q2FYeyGisM+dmNcCj/T3BXa0zM82AgWH2CN7r7RikEP
lDXIUKRqn5eWv3YBT66sCZFJPjBenhlxvRiFwuMsthtvYgLN5Wi2LmOsxA/g9Y+9
Fo6fvsxcTd0m62rjH2/T8LRn/+mxrEqrBTxT0EBZHgpsKeFHxzOh3iNbD9IQ5RK2
LpPjPzQVaXkUMhj5gooM+9WTwjyuU92NezOxgQ0oBPFDgv3mnp2cpti9rdgKsP8H
JEQKvhRgKhv5sm5+4PdXVpn9VFYyL8TqRvFmy5uJbUeL7MH2H4IRQdS58tDvlSZR
NL8ME87G5fiB4d+FYPvGiEZCjm85TJa4lM37QhffBO0oOeFNYyQOyJ0YWFRRD87K
5SBUBwAjZB0VMY/lSOvX5OebW5XEaWVF/KELf11uq80RbjCgYl0d7to1w9IZf2d4
2ALi8irQLKY7lnD8kf/ffvTMLWlFxV/GHaHmdIwDcfE3uijIOZ28ZhEdgLaOr5lp
8+sNJPotKzA/r9e8z9Sidhooa6of7DTFZttdRrhUTrPL4si924za3plHs4TXzP0j
FTb+2KDPsof5RVepIY2cHIxfxFLCYM2iiYSd8axxh5wl6gp10F9sK0ld9IW/543E
tiOSr5OpNyXDp9dQ6jlcJCk1nDDlQwbGMisqMrXmH6YyOOtscFJr0d3NdlEJlQGe
r7uNqDgZqmSZEDv62iy440KT0uyhhvEHuRtNHdzEghFSxYfiYuiR2AyiosrRsn0b
rqF3RQLibS/erjUbV91HOLjXCcQyHG4D+5mLsyA4Vi9Dcfxz8Fovo80s1JTLnLf+
3ogE4QdiJrXTj99ekKMfS5DfDVImRMDHARV4XrO8najeQQtjYXOzLosoMTkokTIY
FAGI2ur/imF/HCVmFM9BILHg9CmD68WoIF2ItjPUVUwSN4UY3dMtDmy7PJk2d5Jx
dP4ViuCEmhiD2LDyH6fsO2a3op4BRVuPBHKCUSdCCj84Av4gZXux5c3FE2ic39FD
iv5d/kRXpxMNHOCLwokOGwSGDmnvomKj1qkDjoW2LAsMWf0DLutKvAIoIwOIc90r
pijDaU9/JRrByhIZUx5GkMFhaQr5nofTz1x/H5pVpOCloc0XlfjLZ/l9oAKeWjp3
qljtcagMI610qu1OxFh0bCQYJSF1pP044VQviHtqP8aLL+N7Qa/SU9WcL4fQU6UW
5FEk+E6V+NjAey6+JcQEy1DWIlXvYAXp7SBCCkBgdCtqo2mOOmzQFIzuaaxvQpBd
Cb2MPUS8aNl93kAB/YYNZC98dDfeozcqOOxVn3dDGxG6XQeYwbm0hgSKfrpd8bV9
na0bBtCTb8yE1nraE73kKRYzJpHCajChGHg06/1ed2P3LTic6n++QIokG/hgDBva
TAKT5DmP8RQsQvHsj+0sSCOHjBkt1aWvMmvOcIJJjrwiaZ6Teh2DN4ubIo7FEJBS
J/QnEmTU3r39rcLEE+mvgUi3C1vssMVC9DK1OqYlojcqrS6K4EDH9P/s1m4aFZYs
ZzhsNzmqks+NyGIyvypnY7V9ah3+lyEXnbPsgEMR5/Vv+3mVYLq8dZvUNfhWQ2/Q
sVp9E1nQc/V3v4XMUcAzFbN4GGVxMH0+GQttmjrspwS+kdF/I5qOYpvYviNvUGOQ
CnelVDXVJtMXQvOV3orXqxBJGnlxSyw1vLKuLkd7Bk7HYEXT81JV/mrEPUTsKsdc
cSwY8/nBlMsaoYf/PzPOApNWOktbu0X2eMR4nq1arJE8lulUq8HfXPL1cLhRAzfc
rkxGl7IYBMCvJSrewd8F9fDItCP/RFpkre81n24rarQIqFO4EtYGnm4/sXjtexJN
GVY6+/o6ec5IJe8t8dC9c0HoTRzmFfQjb0urS+N1UMSYUvVBgVwOU7hepbGf3AM4
g5TqH+eqJ4mGgBJsjd8uHe7noAj3IKsT5JP5JG1iQ/qAjt50M0YDggnjrzw8rICY
HDpTD+IvkwGBVgfdvIMH5BusLqJCVpq8i3WJdzN2/XFCeBN8hWXVfu3r0Aqpre7T
4kpI8RI5obyH0gpJadVYN9elGm8Lt4+DRh66KAW6v1e3cjcwyej4YAG1n+6K0ekF
og8T6Lt01TCigBhTdszOX+IR2uht2TBgKLL6vTabf7EOBN6SqSh756SAQ6ziPSmo
WA7xCKpAO3nnt4wL8uJDOTotKhVrC8kwEWGgWEiuH4mYbKuv0Dvf0pRHeEEa8NnB
8vL1d/X9liBJMuREg8c4lrJYIh5bX9xR7nh6bXXSTZNRJSh/tCSBo9mnNzC/pHHI
/vV9uozvLEgDQPl9rDdg1ITDvA3T+YKZpw3bfET5vh183o1U6gUBMtBbPnAZzRpN
OmtYiRe0fq1zIHnyQQHEcwYW2KOlJbppRAON614CGlPSpKdM8uoDW0kG2SWyGXAV
DM0ljpCmJN9vvpADsHCAE+jX6RPspHxJN9RS1LxkH0gadpLtNi5vQP9NN9mtuUgE
hG3ShEs1ksgAS2lvqoAKUtCYTFTjXXg1mQ40mmAL7ApdsIpdCK5IWiDj4JiNG3GU
0mtUs8x3fiB/B22P0J4ZqtVO66heR1CGal0EdFYEL/4DXBQ6M0X4m2MpRyfTIH1U
S5qHxz1h65r3GbzU52qOLkLPy/y0MHlVBrT/eemA8HY/cj9Zs9gPXzVusnpQAp3X
U64nqg6d0YfatcNEC2nNwXVizuxVgNMN63wDWt9wIDpZ/51I6aEidR8Wg/hLStjC
ffoFYn4RZXuaBzt7M4AHBc1t79fSUKx55l4sxue6+wmmSjXqVnYqbcyFq2V5ycb/
WMkHIfD/g+hJIKtCFON415UHTYHaw7bX4uj5dC6slH5OrXKStrNh3gv5oTOfJkkR
PrCwznnTuCt5SwUOVKXg9nGh5dyJvCxwLueFigVcY7S3vvwN/nnoWS2fMFvTn7WH
1gJ0lbGJf1R5x3Xi6Lgvk+txKwoKeFFxP7ZxmYBr3aHu1YBtCsSZOAJ0XGlFdTwg
aIYDd2UChjSU4V0tuwSXbJ5JjQVpome60QGxvZrlJKH3O9Rwwoch7Zevnivz8tDh
+v+tNAQ+ak4wHGKFfxNxPPArZ+yqXGJl2Dpjt3pA4K6epyvCuZKZRtx0i+maZCzR
SOVSvyBemCLZAcEnm2kprAhPGQAKk9NLB4ZQTb8ubR+I/OBnr1hL4mUiFwdq1FDO
YXiA0+UM7FmvxCsNqHePboXn6jIkiPwWA/eaKiupEDV06XH2zoajnNhmlMHDHV1v
E07XhJV8o382fwj+VZsCItSSUD0EErDUgXjF17Qg2i5OgW6ox92t85rz1B+cCnME
n/L1C1MJrudWAsmDV0duz0Ww1woyEQp6z1S4RnorTvnI6pJaPCo6uXsSDdUNUrv4
4EuB9wOOzGstgSr2EV+WtNz1AGbARO6xmbwZQK8o6n4q2dmzGFXnc3NeEJKfqCX+
KrQNG6Lrdlvj/akknQuRTecgTA85fW/0q5rKg0UoMjV+kcYWzXjuyURfkduQCmxk
ZPCAqv8znK8P3ygAJnzriwtx7D0DnZe8ettE63JV/tEIDxe7y3N65lXGkhQcG1O8
cAN828LftEEf8VZf2l+xtEjfqO4qvE9SprNtJkzmRVuTXxDInHLYTEp/Zdg5e0Ix
KBdOdOd5f2czX12HPS2ulv674bC282nf0yh82c8gkeQXZPgJ2RrTFBj5YPzLnwwb
lKw2E/fdMRkB1HdMk0Exzg0T+DTmsOESX92CNKATDINxsMPvG8xY1iTTTLp4SEKS
Y3bRTDFLGcjWFXbUywONiNBRUeYNgui0XzIQdAPHSIbifD3UhmiLezFaMHtoELNq
HzxIKIC8MY7j/uwMYIWvOuc03RpNz1n1SvQ5ok94qoWKGlAmcxurfQhfs0TGGxON
MkWxnBdDBiS/hxF9zdPf6f5G6wXORL+sh3PU4dLflyUyvvDQMeNU1zkZ5b/ElOqy
eTz/dgySRRqb5zdxQcbmR1OJJPG92Q82TsuuU7SaLXisx7niQ1OEapo2SObI00Zv
gaWAe2+jvml3aB3aGiCKL4ZEjqso3l0V+7Y+Fa5ylrsoUpyI57uW7rdM6317VY2M
MgD++SxNQctYo31m1qjfpezdT5/kNjbNoanaev/HLoEqQlQq9Jri83qFDiVSn0JJ
fxzxdeu9SzWKKdOg62YxN8t30MasrOsaKbxW/SO4S67DtFGFsEBWZOc1Ie5Gfpy4
EEWgLO63zsXfEpha+KVxmJBx51WYJdR3lQGvOW6nqcdE/yYKv4Ec09cahpo4Gs9S
dfo7EJNntMi+odOEqlLM4H8qn3bM7PiFD4pF+CLtknaYybMxHGiaxYzTeRzquNWu
`pragma protect end_protected

`endif // `ifndef _VF_AXI_ENV_SV_


