//----------------------------------------------------------------------
/**
 * @file vf_axi_slv_resp_cb.sv
 * @brief Defines VF AXI slave responder callback class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_SLV_RESP_CB_SV_
`define _VF_AXI_SLV_RESP_CB_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
q8jhzSzURlQMGyJULS98jUikENao8fegXevs+IwUKbwJaRLlxoAHX2HPtjBSHc1C
xNlW9vuJuM3lfhgKzojEiUJloZICUgP2HPFCOQFKEw080mZyUHIOyyDGPWMm1JHr
db5QwRJZYlByKevv9ICo9SLmW5qYL2NyEtpv9v5rREHdHbR58gHL4pKcWCEH5RWL
6HLwO9laUORw492yUmREM8TRZRlg84y6HdNfofKrCOk36AqDT5jrRoo4JPK33Ny/
2wT+LoRYH1tL4+GE9o7OnAGTM99DhDCXRmFoVTEq+ynQaVuoyz1EdcOl7uAuzMDc
coyf256qmdbUCrAObcI4oA==
`pragma protect data_block
t8CWGVB194WW0oQQPQxsWqSyZ99VzG8SpXLzb0E+19bQTCxqDZ1qOQlrZCmOAFel
YvbRAtl2HF52pgQ3NKa8J0Aj8j3/n7y72h7QvLlSHxtqiPBIV2EWlE18JteubPAv
h0oqg5SyTyMD5LQWOed3dphDvAZkImsc3pAWQnX/n1bm5MHKEkA2U9dMzowoqTEP
wauq3BcJd3i5ILkDfW9ZXr614PTF+u5FLeoLhneb/DjCXs/CH4mLDIxwpT7B62p8
7X38p1S+N9LcwF5TDBC/GXOcd7+p2PdAf/SyLHhvExvkFYPNbf9fg9Wh2pyvjoV6
bvvLxb55qebgolX4bmiEPDLKXM090DdFMXy+IhqTRUBH6Ih04U8xoE8w03qtTMP/
YZThdeV+2oMeJDlfh2j9Rns5evRUO6w22PjR75/ISQ+tIeh8UdaZiq+xZQoWSg8x
pNPSJc9tQPQLcbw+lYNPUnhrmPfX4H+IE62GkRAdHCWhYTf6Ruywg/hMVCF34Np2
nUNRCY63RPut3g+jWERUkKVKWtcDGy/GHienK2QvtaZpk8JPPGOZup9ppUj7g+vy
t9fFHSQvL1V7+CEuvCFjtZO0zeyV4Fd2FrlySh/ZM6VXbxc04Dv39B31/RwCMa55
kOCDuEmi9F+WKwuSnb59GmvaOnFeq5FWkaVF9Yv9zMVqQ+nINWuwDiNciV7kTGuR
XqGb1sdG6gv0iF7golmf9az9gOmXqUtVwa3KfbTlaAbwyTwRxzfLiVADaYtFMLaS
omNS8DcPWwxI9sF5dyhfk5uK+RL8yj2Ej5ukv1sTs7fv+xJnsTE55W4VZnJbos0I
WwrBIq5f7kwkMIRVqW52GsDfORQDcYZ0r1sNaDLmTkNjj5fOgEyBTgMBKY1spPqb
W5C/QN/OqqFnMWSH4pEW8v7bNtCFP5Xm09egSMVk++JxQQ/Yp5r93QyDCqFCV/Uq
/sw0GvlgI+aQYka62Ukson64kWK5R8pGl7wY0KTtldjGfnrfd0WZVDRhl97iqPIt
lGKKZ50X4IN1Ay5m5d3kIX3pq0mh9GrkBu1z2/OzDqzOs2h1MKo5qIO11ye9rg8V
EQR8Xp5hA58CW04UccjY/4a9Kfe790WqvM1IH4EUrBsBKYJlEHQLWCaKfUjyTu1e
tqi2fn43Ib7UM7m79Pym3bzk7Zz1m//d4ia6IDLus/D80anNyQX3yJRTkdmSdX2M
syafc7500qA154d1v+X+H0ZG2ZNYo6VGZyFaHRrX/9FH/aQBXJChIsAa9ZJArjnE
hSneQdNTINBevt0+UeB/0EMbM2MyXLJgk5wesxF3NVxNSRN9qaLvu4uX3MvufRiQ
ViAIgCwV/yVftOkPJ7xMdNw2mEWBVeBJ4+faJY8ki0+lQ3sucdd2c7yMUNikYpxO
8xZEsd+AKRclnxI20eBW8ays9dq0BsIoptdw5wm2P+fqeTtkBBUfuiPO+kASaPZw
GKXBvBWPGG6eidUJ5N9/eEpQYNjLJyuvwXX5ChPKtq6X/l3aMjtNRk3IhWiOw+sw
1agDg5mUGVINMuQg0s2yQFycV4+08Xc8TtooxZj0Ourg8BjMFURqosvv2O2FscVL
/5C6rffanstqQaA6neSdk4qMqcfNaTqTsUV55JuKtG7d+z2N2X78VcnV2ZJCCdzw
LJhVRBxV0JXnCdOCGt4HStVUVisfGL6xWH0yX9tJd8X3dSIqiOS9U21kicTueqmS
P7RTETHwe/Fq4Xeg6QPL2OFvtCDbaETCjunzyKB74OMt+BAeD32QYATKhAhMjEui
GdV50u05Xvx0FAxyOwAf5DCWl4A4rXXpolGJ4dAkiILhYLv5ZrsijBXCu2K5yzpp
HvppU7EXk0mE4cqpAZSHsM+eC6SLya9H4pmPPrc4xniRaocADIL0ThOr2q8bwAt6
VCR+6RSUmQPeFholL60ueZCeB6FPv5j+kFcBQx4kohPMceLKUBflHrF8kUSAeiaq
jXavV8Jjww2HFU4Qcc89CPFjnf4Qw7+dPw9P2JYXztoRjxGs7EHSq3on8uGWwQ9Y
Z+UoGnstjjgfY7RrGHpabea21dDSnchzAutmES4jdpUCEpeF+6Ic0bV9f1Pjc8va
1kEwBgfQBlFLJcT3rI0hXd2FF8BTJndRCGfeDkBr0IeYnuDoN5jwtBOYzZrn+0re
hijjo1ImgdmIwIo8guj8bCFulQlbxgM3p2P3fyRrJNIKwR2ibxcycQYv3RbpSEGs
+eD44A4rkDQZRDn/yNEVHFoQx12TTbZULIqJ9tiCpGvL3di+Wl4dMtmrP5+mlOY8
/QtUgVrkbFLD2t9VsQtF9YicHtBX1SAdqpF52R6sUAQzGNy2fK/aF/q/QnzGfoea
uX93YM5GFtyfv/3FOEe1zC2Tu7QVFox38RijkoGnhh1Un8LHKlVCT86SzECaPFks
df2bDRRtaoluGSfddckQfGPChrDm0UJagUO4mo6pbl4zU83CDacHH1zmsZsbIyQo
thEWFkKJdPKNC26n3/pCNrXTGhRmSZS296P4EN063yHO76NcouO9XW7qVdrlde+I
TMdFgTcVGkPAf3NRzF0y/RvrZGbxRa0AvlrXcycvLwSkIR3Xp4wJKP0UOv3E6WAe
xHUnj8UhXQLFK+x6189t3K4kyWW09nyT7HjZg5g160KZo3HkhFyPjBwbICrdtxP9
gLIr4YBdajt2+9p9TRR68j5ksVXRcHMraYgzQ/XKDwMbx/183eWcvlI8/ZDaXSNq
NiSxGbDiG1j9tTK9nJM0Ahl4q2LsanuC1NLOfkbPUZQuzVrZvLEOwXXKYxCBtA/x
oWvyHE9LJw4xPPAN7gU4lo51QxtnmBn6x9cIenBne3qAZSHrFnDCRYzYwImiIUx/
PGRftgV4W1/WuIO7K0XU7p7sZdTaug5sbA95PtOLULjBlCO5VbccCteeWkHOVSGl
OsTHgUL39AsDQh1XpZEUkwyB1AtZghRVyzQlzE6fI4ilzDP2eVDti4SL1PWG96xS
VlT0CFyHhvyQG8tqFbFihwSuX9O8IQMoaaMJjIXjqL3WX6o4oN7IM9x94RFOMZQF
FmOW407Z57atyKpXDUKhamKwefcYT0Yj2IBKMsfDg0c1jAwt8m1aciAVEEuEtSbn
h2Y9gFo/8SJE6rDc2EvIF1SGePb/fG51qbeh4oWSSQJT+smaCq9y25zMe3xrPgdi
g43r4Zwc4ooYHnIAR4c5S9pH0vEKwzxqzIvFELyYs9yVlrusSGtfmm5SSSaWX8M+
CKEBTTNNCCLxY/3eq+DQpHh0T3wOhTT6NpGODew1ywn18q3+tHAsQSB11PS9pHHV
BaGQE1CUtD8jK67VS1WccdBLeKLVSU0VK6nQU3l/jXUWv+MsGcWHqe88KBfpPVfc
2pyaYgua+lGTuMLFax0IFYdZ1yBHaNI7IVLtXDD2GNSNlw7k5kdfPuQmiwxHg+/s
ZMZR7/TWJMLNFQq/Bhn7JThHzKdcVz1xALYbgnsgq1C6NyK/BKGkYRDT+f9vqrZF
xV26+ME60z+7lt9B/JP7EDD4M2loJKTzTv5fY8IRUUSeu4hfT4lN48ddB0dP6esd
6UHh4CcbJL4ApTm+mIEWL5ttngGah+Fn38+va8xAOtPaEb+ZfopoYi/qOvf1JGkY
liflXzN4G+UkoT9oCBBo7tm6lKkJoMLFGi4z4fClGrKSIdrjFIjH9l65XEVRMmgh
tHiPfqxJhzuhZLTckVtq5fn9mkYv3UTdsTjohd6V3KEBmQOcMoKGbGj4nCng2Qnv
rVDvDmsX7FnEd9nYX6sqegoyJjGIvHVaVX7rUaUUCUmz6Y4Yki2nJisdG5qCNtL7
7cvJH9KUUd4UMyQfKM+/pjiShGx1WzlRtJ6996HBYGana6tTOSIjZpunmoOkFwqL
kGablnDe+07s5xPpZbq4Tkp0yQFEQ9fEq+uPQ4EtA7bcaeNPaLPfP4mXDjOdY/dV
ML+enLJjuq4LDOBxJssJwox9pDYyKwA1OHQAoOFxjxKgOrwpytoODr3DYIkkVxaa
54qustn5ZUJXEd/MGzBlO7tEfskmu6LPMSP3oO7A3GyWHK9Ud5U6UjsM2K35BLIu
fn2zNiwIXFONH0OrSxTDpc+72f/I/WEojScRDggW1mbHPaeQ9xO3X87x4uiP8/X3
RhcN0iceRntIaQfNPRASN/tQdSsqn+z9bo+TPmJHYJOZXyRssEoyNNBxj0IyaHL0
XpQbdOK0qKaYOHn+YkmVtZTJABl7Jd+Sy4O8MX7hZfZa3VeTbljHxSTC9wpzXOE1
+37+r4wHOcP9yM8z6xXoT5WCNikm3KgEQioGxb8MV1dm6f4aDCH+ffkCWDwtgcGm
Q6qdT5kwKeRJyLPLc3XTaFkF+xKoZ0fNTcOr+/BzgHso3KmE5CVTupq6c0hhfi1s
yGyvlnslyj4yQtu0sai4zDBKVsXU4qBH/+UzIKDKBj94iavjTjHIQGZkVQ/jtuSD
DfP0JbcUCd6RuMITpuifLYe7tpxe3H/645qDu2cSr2R/SsqW0veypCzSZa8fuyAN
ct4ylPRaG/Pkj9hYksgCIc8E1bLSHUa4E6cW3AVhd/Lvlv4A8fpk8hSxzE7LShaw
gkbZ2zrHvXjXYC3jGuAfPZ801ZfIGg3F7TeTE2dOcPbbnMG4uXq5cVAUCXE4Pw8i
rYzz9QvQeDejDauQlPsshZr/bWmBJ9BfPKfq83QG2DCjm8QFTtGgHodfGS8PF1pn
OeHmOjw9FOdRM82WsKTKaKZmIFgAKChYa7lVRIkvPlwzLIVNaw96GSkEWiLtY9yc
PQBb2QO5OZ/W7QvHaOxX+b10sXM1dgX5vivmnnre+pFOEdq+TJ7j67NDYZc5IYbb
5Q1Mo8k2w9bhQKrPMPaY8vexIuzI6ig0DO1dAT22L9v+iB9rgjZglkMNWkvXC4bt
xzpPXz6+TL/YBwxa4zi0RhLoA8ayaw4mOHlj+EencV3pL3BqNyuguO0f8860Iwcc
9XaSkK0nw5VbuHoSs2p0CoGyAclxl1hLFbP1y5GVPx27o4fmQCzWLDV40YJQGwhe
Hmy1KeDyn/woSqum8dHwmyf0BP0wBrreVnjKRaRP/Txmvy17VHnwyGeny51PZgbP
QmQbuub+X3cmMtBkwJlfSXzSFkHIvWdaMh8CQRB2vl2/F3rcUZNnp4+DjyBl/A0U
1NGl3TfgUxNf+LD7flmDEE58tcl/7LHf+momPvEgmhNOH6eVhpaBwxklIrdTrMX+
XFRt8OgojauTL53ALz2LhICbTax3ImDfRIjd23deqgQGxGw5OIID43uJjGCviyqp
Ip0Sy9Gkpz9mm5EKFvXWOFmT6Z3coNholPS8epM9G4KHDpobwlzktocE61V2mpeK
4Ish82cjJp9zrTukKHGo4rjK/IFKX/wNOHCE6/9koXV/Ko/uW+L8IYGriWx3a0aY
XW3A60q+b8zctGXHv3DhB25GLWIeSTD/7awXFUxAR47tDhSYCyn0LsKj8YhNBJ8L
TBlkaum0XlYSKwZc2bgy7LALpaFT4AykvGIwi6u0UrPDrHvHKcRIo2EwAgW9VAQe
sXQ3ThvNIHb2rae1OpOGsyWIX2p0JaiOykuOPEGg1wUmYvv6vYV6TN9d27xvPjeM
dZkgmSkhH9QwvZqzAhJ6Tnr4T4xz23q0LJ9Ho6p3QwxWgA/d+hOZOxJj4nQmP7Lp
IK1OLmICkYfJs2l3fVdqPWG1FnQZ/KS4vOjjRebh3ojB70Gd7OPAdmAS4WG6B7j4
D1lJkIoGVt6nV7FP3X9cnAF74vomwhrPLZ0uK+LeP9Kz0LLQJdkCO7YiluRSTVUA
Gfsw8PQ5UMxTwUW4RZLjsHCZQKrXvhyj1I2tv6lrldUXGPg9+5660GwNvvkWM7yu
mGQrvLqLmhyfQYjBZNzJsaqNljrN3139xgGN4gnPdgHFb4++79/iUZdwyt5URUlG
IWDeAT8JCeW92Hq4hi5gfKyHWtSFHcU8saWQeOljhOkC7PA1JAtyczuZ/kT+1AqZ
hjgYfVZRZHJDQd/DwcL1m2x6PlCIYLflBzF4TUXfkBsw2z9cMeSVVbYK9CQ5EPxe
GEQ1irQqYe606mEHCF/LzB6khINkLHW2nWqhfAr+YuDwEFhrio0edgB5DB4+f5VS
XibNsbzYbn6K9Gbs6ZK5sfLur6kf5JeqPHv3Aju2q6IkksRjRD/9W5k2pnPTRZGF
6B02UdJFg597VdeewaI6JIOyX2aqXxeoSfhHQUXYu0CAXddBjHjwUwNTXmjeT10g
iEM7z9ZF/suwsc/xFWH7tc8L+t8NJCTkXnUXZsQ0EdiupcEpzX2mwesaAS/9fOAn
kb9R6nHMmfGoUyPlGiYGGfMX4evU1fIRf0CafIJe596uBlNqPhx8TdgU9AU85zC5
DE56ngvs4RdeCjjqH2+NHjxwE88Vkv67hpJa3dgTumLMIiObVYlMOErCHHfYgTaF
BTbuqaA9RDZavgXar8mgt+1j7zZkeBu7YO/v90xeygbtwVZ3FodMSXE4viQc1oA0
R/1uvHdqBpP9owtCMzGsP7xnP4dJqukU4nzp5//tB7MRPkJYqRlbud/zu0qGvpSa
1G4Z9W6u28wDKitoQwQJ5ary0cKcqedyorGE9AZwpLKDGZJ++UGSGCfUbeRMwLgP
/7YtMQ1WHHO73qwBDscuoh0Ks3Iprhw+xoGrh9d4kMI8v7DNPU46QSCOyxTtWfcK
CSsJ9Ews2/ZLc21hqOrGqCjzX4kLTUSRmM+Zp62xxGQcPCe1JPLmbXKc207r38yY
8xYLoE19XFR+bwMYZif03hQFY0y8OyLHc55jsReW7ziJfhKUKA9izyV2iN8cObUZ
JcfF76tNTpIpCEtztaJFO8ERervbYVHZY1bR2TNZ//Y5fNF/4IT3+UFPG/h1RrtT
bdXZ4bPgL1E8F39pdnJ3VcovF586lcCE0vOTe/vDsohaPvwiU6I7Ej5xrTYg5KYH
wCjznI4z1PqnHh9Uve1helghzSto2+D5fR/ElJO3pm9j++UkrxdF40cc+SAJNBr6
9h/UK+j4hdLCtDdpl08MSZg9cqiQZuPM8CkLwo++5c+Pr9bcP/sHMOKI9Tv2OK1Q
zwh4yx8Gy7MgBL2AnszTqmp5+JzoaB8Xw/eSsZy4sFBscs5BWve6QvSYPJR6HFz/
QyliIBmvK2tLKlNBfywe7oAFevJeY3Z0dFvdtnmhgvSrc43nILZNm7fSYsHeARg6
FGYuhXihlvy+v2uDnX/9wS15Rijwl56DbsjfA7hXjn+VF4m67J6wWreUPMM90elz
4BUrK0mFPxdtdBQTdFDaNkmDxv5huKp7cT5mLaAypYmJvrdrp1P8a3DErPsbyTz2
CD1pcKG5mws8AKkaYXnHVJCfe516/GWFIxktbR3pBsWrl4+lYPjUjcB3wQKDpH1u
e8bdH/z6s7H3rsSGZnVsSwL5VwcRyeK4E31/mOHxb2v8GyMRgoFHODp28dSGPDCd
1fdsHh/n/wAv+hWUSp3SCBebmTJQPQH0dnaJ3q95HVkFP8bGf6hJJR3YTNYJ9v4c
3t6Ljwp/VSpdsjKavPQQ8LCaqTTuTCsXSY5ehuGgvCocCkud/fAwvkyl5Rjn9VkU
Pd6AWs3BUkpB95a7zini6/PWrE8cjOvuwAmrwIGfTCG283m4tPgbhbzcInFJQ9zD
OC2mr6qSrsQEJmal/03nXjAZ6wl/QpuRb1hNJZU6H0+I/GDa10LsvxRJL/7JgYsP
bg1t51lka3h9T35FIUxi1zEaAEVBnTky/iBH7CAzLnxQpS699u5zJG9WMtFFi+bR
lD12yWcAnDNWG3hp1XhMf/hI7m0zy9hXZO+o7U55IQjcMcCmGkHbzBk0HPGhnZir
UlO3uJE6yzSZxjNht/iFtAVmZdqB0/w9NsLUNZzIfh6q74DPOVZj3CPkEs0Qhe6f
mcWF0oQukARQ7j2u+KZyEfQuHJYjBFlxaonJCkmlPyyF1h9aipc2TiOQItnEk49j
UoMnzwN/71FU7OrgtRe9gmI1hAs+4fXJJg679ymA+0/rPblv3x9cK0ctSfd4qiI0
wOHrd5m1mvD3/9w2VPckR6NIExPsxokYUMLKdp5hYqnKGo9dEtkwZyZ4rxI4vlzU
h2kv1iREFSth9ARBG7nT5AuVSzA04fzl+SD0d6iwcaAUTXx6gOnv2PY+PYyUoxKQ
DrYuF5n9D8NIfschO6T2EP/ybzqsiHVGL+s68oZhArh47glw7iEAch9FOpnm0Pfq
Id+xN0gY2pNMJR6OtkE0aHpgqdPoT6ASoWHJ55f/uTwJf3ExR/i2m+oxGVW+sUUl
6ZBaIOWsfz6sgixuiTiZ6Y3gfbeohn2IQUGV3XRoca0DxxjfFAUDm1lHE4JbSQVX
M10XnUqcLtc3bB8eynSxL8HsArdV8JK6N9fO6XnswuQAJ0xUQ80JGH3y+Uh5Xf5y
CtThP+StNJzSuE12jbfVktVjH0zZ7VLdf5+JRkntCwPJmKKQcDLvNIgSzzqFUMPy
IhaCYeduL1JlYpF6saBDmeNSNcOB2/xuv2IhU0CBJiKHcQZ9HKZNzUfzcjf4cYlt
LNup2ARfI1moXMzTzRfpUHtUFYKF+kYSNTE0X24lAdQoXErOPCovy+XL2FCcaJQY
w/l/y0cNirje7B76VXhEZ9qxMeYZJwmmHEK0M0BO15HvBIeLSn9HQMaeofbYil7Y
kiqDX3ACy9w7xpQrrOCAywrY1yHN2dbZDH5inCpq/e9fBFyy1ac24BKawBM4clkt
MUmB+3L6uzduNfnim5BC6TZ1Cmeyj0AUUvo05p/yZzg16/R/Zlr9Anaf0oup2Ur8
MKTU9pW0bZ54i7a1UYBBwOKzmFRdpna9+lheBxq4RMW5aySWtIkQe96Kmy9EQ4L/
EnkWdkcmGyrhvqPrHSR+hJ4Evw/lwzKUs6LfnMoHtyo2yYC3PjxXsxEkZOf4vE7E
P9ONOX13keB81SziDGMjsCpgIG3wP4rREN9+dg6PGQjVXxS+8hUNoZZ4kuKmzTj8
hUKgW4IBomB4B11FK9LRkE/75CAJ4XI+YG0vRbw4W62HucA6EDEXMxl53qRz3DYv
q0+KviZkE5WzobQ99IHocVp7DAs58m7/lYSq6TrKJzpv8AeHPMxsb+sOQXMczkWD
oyUdAegPJ83o9frGKuTG5aQmBH8MY7DWkNIyWFiwfQf8UKHbi85so3FfOlawADSI
wS1CB53mu6HHwmciHkR2IlwjvqkZY60obYRU/aErt6Iif6pk2kgYMQbgAjH9rUGY
0M/i5X3alg6XfLg2UXaYIDL75yBvQBJ+sOCeJ3DKOC5/1ZXSgOHjB7tHzymBU1DC
VrsoY0twetqk64sS+G9MJ8iYOH7B4JyIzaGsH+3RU51X4RSl+17P6I3KnYcHaJbN
9x1fyhY1RxG8DdBjqJjaerGwPaZJelCqT2uNI9dSXqVhBhxo+Ohwhq95HmsMkiqW
J1wa906QdjLLbe9ck0hQR7pVdBlloX69Cf5npi+i7xvwBitUk4Xey4/EIgP8Sfig
0qrHihR6VtSTn0JM1d6KvReWfbRBOVNDmous+gpa50hVgUgtlXLUbpNe79pv1hQg
Y40bXtvCwv2rYgfq3SyWci5ZMav3YiiJrREpxAyanx13PQ/ap/IMf56X4emoPp/m
MxDndVTO5hr/5cn7I2Q9t7Mn86uil0P7A8z8UkdKSA1ImFWa4+GOMNwRH1p739VL
1ZERY7dzHUEFgmSPGf2Tv1CMCydVmIhXes9eJdi5y3n2qmAK3FIgcfD9jG34n4q3
ZY9G/Vpf6iMVKlH5hNnoxsMZY9adcTQBM90NauTs7xsdiYvX0oFd+XuGQDtDib2i
y8zhpUO5idOmEp+WE/j0NuA7096GAfXxq/PoM6P51N9GRsrOGTdipPfqPGmbKi2W
cwRmJApaZokNHMMWibqNv90Z6gsofUM/uA13/WFdt6twvRP3UPfqTkD0TNPTI9/b
pxPlJs4TPRPnJ4ZYfKBX0q+O9Nhki6iazvIaawTrGIF23YVnOPRQrldWOffgZict
NEBKS6WEb90/fT4Gqg93fUDSyf2Jt5H7/grrScQAsqzHkJjjawWwC5yjavIXjYNY
m4B6R9Xs36pMNipkmogpnF6FqgUbgaQonHGL43gOO3a2nGKAI4j4JxS/Pdbf6r9w
bO4QeQgCK1R1wqgx6JPES1hiPucrYW+M5zCWfjbo1/E6k/MhKh8C6CplfgAGBXqw
jKCBaHhO9pu51KxWSw9MMrX3xG73xMzmhxF6BQV1i+4PBhhoKH9CGT0IqIuvOfcf
aKRXhV0DcADSDYXbixrzKHK2Mpjy9CLk5VUTtA7GZFwxCSpcWhs+37ECoxdHhiNC
8B/cuw4fdKmSoA7qYhW2XiG3KrLH2qRCqu56+jtVAstZQUBGEuBQrMz5/DaCWY/+
uJn2gAs+0pTGKxUXzXvq0PMNfWQ2p7gbJqYkkt9hj/Ntkcl8Z7npQMttaoOCM8MM
lppwgXSLLlFf+xcdR7pmwYDlU9T0Dy+xjdO5HRL919WJFFmjBzqZstsIUdGuVMQo
HOH+5mFNbVHE+tI1s/aaKHz3p1A6/crmc0ENUvO5kPvLK4XUzGteWr2AU89O23Lx
CbnwNmu2l5+lVj/FvXGaf6o9AG39gtxtjkJOLghFtwdJte3dB5bnr86z78F9YG7C
vh8e4X+TtN3wwvPLiLmo9j17O6SWG/lOJKqbl0/epIq+jQCiDJN517SxWv5hfTyn
l2MXj/v0E+QoJ6ub2nGnEj44MtPbcNsNgH9foE7Z//Fe8EDa38rCKRPfXiAmIl/o
/okoFL79UaYog6OwQSd6yjhOJtWuDW0xVAxZWTqpgl0jfo3CX2d1CGfKr41j1sui
Fi9GthOWo5GQhZ+nsdhB4Gu8J7hsEfB0W/Fw44KSi31hZFt/eE29VLInSUh7uSK6
fX31NfQDKwxi8w/Ig/+Enohq8iMjKA4YJHcPerWLcl+G9mrD0u3X09JmjT45hD7N
ikyKDcU1l3F+7HEb7VuiFQXUzEvj45gNYUO5M0Z40+LTf5X716IswHKfAcOAR/pm
0Em4qmClhRvabtvadIU3xfSVQ0ez+cqm7QGIzrVZamLBySUsEzLXcnB4CYEeksZl
Au9f8FemJj0Y2Ol+OirYf17ZQMRk9D8T4fi5GmhbpgvqIuJjBtOvA5msc4o/6IjX
1JuB1PBw+f6sZ/gCeNJRI/kjrE5FB2VZ/fa4eNnW002FIHQ8aEilv3lEq0QLPAVZ
UqoaQOmOCYLKlK9XHYEEWipponLIQ9/w4/eGWz7+B5zxnyUJvWxjRqmw+wvUP+t/
ajEaQny+Em5SkWTyHKPMPCXCw/S0a9NNFJEfibgX1k86Nh3/BF3OYLZUBnonO02D
S1B2YbdByV0CvgTmY2BXe8KzaCFGKzQs50Z1FFZUeTVYmHIRFz6DdY12zE4KkMX1
8+gBiYpeB72IhFppmac4nOD+gMn/Jnr5lHgpxdJ3ndXy32/4EN2yofDTe32GdLxe
U06ro5BeQ7UPD0zzOB225jcZaoo4Eh0ChokaF1fi7Ebur5pdCfY0ZmiXZPgIsKaq
u5auG6aCuodx/PogYOkK5PB3XQ4P7A+73bOtPMSHhK8wQYE7HtviPDd0pmxFNRCO
Z39ZJLrrODRrzeZOsTkdReAi7GMVf0cFXYUV1Fr0VKGUxkkRoiP26/cWvVrtdSxn
B//U6XMeQ2rejCE6fyRS8jKqbIpTp0EMHpOZ0ur58nNnOQ8hlTBnJtFWHgJoBj7p
MP7aiHRmnT6EXQwOsyJLg0DyGo8esxxfdNecrJFYn06Hs13BOKDl4Eis8MAiWF3B
vDNDpBhpIOEbbOK9tsGy6Nxea8M3dXw/uUMfUZswEskesUNLEW0XMLoVlmQv7udd
lPb4tXfskIsw+ZoNP+kHZVtjlFetBlCYEk+4WTsotILfUxe31KKE3o0IMUvKjPgY
0ibudh1bN/tdehv5XVmF81eMiX8TtHmmLp/l0IcnP6gAD1KdicokgUNoIquTOMdI
R8e/u6Q6inwsFM3MIjAGKTjnQkEGsd2hOzBDfnauQqas+0LWJXMY0x62/YG/NSa6
1yzzHscrzPhdX0B9u2sqa1e4QloAuGnxzCTfScfv3MGudZl8j4Rfu3G3gGNRggvP
jckXGumTxxgn2vNPDPoMaVFA5gEdkcPyrvAqHNqagk3IaNuFD75NJCgk/Fkk3Nfg
P25nuYfOalCUCqqZ5i45sYjCEw/tSVKVuCpAQLRVymBae1o8Z6OTiy7pLTtgpL9T
DpPb3qcdxebBmy2IfrBh7p6gBgRMT6cx8mOe33YWC+cDNaw6pHleRHDNAx7si/Kv
u2BiD88hpM6jUhRa2Q3iU+uVyqwxR+1pRyXcX805N7I5jgcSti7cJLtr7Thi3ETA
RSpLVm/Dxq6c58ocEmafRUie0GEMs63pXXbhrHJZrBgcLSF+giVR/rJt9FVVhP2a
sqn7fs4jJ+Y3kMWZFlv3lEHPuwaY95CQ6lK+jP8tPvUvAsqDhsC/lQrsEWB9bPw1
1R01Cot/9Efdm1q8NIlb0lKMpk0MuZTkjAl1ftj/KM5zuhehmnHZ+03aRg1chL1V
2EqNvUGa0SD/j29XYKf9rsuQLq+n1isxdqf8r7/ARiO+iYSdfVI4PW2qbiXk1sOr
pUgEGKc2moFMRJrKucRG5Ag58N6KM82ro4cwTCJab+dG82gqgfNLBFsvSe66Rnz/
RmknUf3O7EkJE9U7bpN9aYNTEnNaW1+SUNaZLIM1nayIXuvp8X9ZOJAqO7jXt/XG
uyj3yP/9H1Yt/OtKafE1FU22NNBzZ9JsWeuqxp+78LbpbKSMX3b4MlBcUHETg3LL
FthaJ2o1YzXfUieiw0WCb+ylGO9zTdDIP/CQIEwD3W8XRfzJ1n2itohHAiivjAc0
82ISiZSA/66lLUh9/YAQ2aMLv5pLS8cvYeFzA5pHHaVsYFC5O5mjpxwckUrf4vDN
DGgfMPOxKW7LqUnC3ElqDo0nKbilFnl0imK4bh3YywfMvQIW60L8knRkNhis92xr
7JFhNLgwU+JLULCi/bhv12GKhr5urQejO1Oo4ucfZtz39rCU3r/2QCPkh1olP5TA
nNse3bsK7BfdLoPt3LiKdCaZj07HrZ08C8qnZ7yWUIA7rwEyCiQwH4oMmX8taMB0
TxZzTjbhpKctzwR+h9geQ52OmIu86fjDBractzQ1YLHPw4j1AeQUng3iAb7LGa2c
VFnxGOELP5TVuqPOsunbrMgujR0Wx5uTc1/dbBjTvxwBF9911mR7zplz3PXRqEe9
xceVXPDy0Iyz4iDzVfAbXgWSo19aVPFFMDld6hw/lIp0iqTQIN69cwdogPRYGZ+S
5Ocq7iUnXCMovrKUCodzVb9dROrNcaH6VcebpOnmGhftU9+If3RKq0Lf9+aiKVVf
ruxXedKHzYtLhgC2lfOHHmIueovG7OEKxyTjeH33I2ogKuwC+6/LhGULTUQ1r6an
5QLkpBHCAGB1MDCJQK7K7vyD+ejlDlYC4QZkxlMr8xgvhOHMPDIYjWb+Ug23GMRe
wd6mDI9eDrIoND+jB37hpQAfKLwGtuc6o7LxKZB4g9w3SMqPkLqLvs013jBxmCZ7
q6af50cWhtkO7jsm0jIA6YVE1pFHAU773Qz/r+bZ/+pc5t8qhS0OMFwQXdDCPBtB
gPY+g6MHxdxlGR2DevBt3dSPJ10C9G9+yWWNr6hEfDhOgyQ34nNVGDbAdkNpIE8H
40+x+DTvmpom90TL17HcMPx2u4Nd8ifzcb0FV14CluaEOLgL/klZEtDlYRiq9zZv
vg0KtwvA31DnxWrXLLtURiratZTRmi1AdD5RZSafohutcKx3VsYxW4OgEdPZBTBn
tm+zcM09C2HG79nwnoj9i4WJnwO+yDz6sGKFwmwwE68LGbDbZYhFoX0Q/IOXy8fg
qkY8NdBS68WVGsKjKEOumjIoM8snB+Rhz/7MPqYw04bKprnkve69iTBq08xuNKmE
EhzPeijG6oXiC4tC8vNLsFeIwV5j6CSAqjm3BqdbOVB7ECZ3MxDO6I+j0DZCiHQ1
S4PyVApJQL+5d7Oh0EM/y4pfTriHYRbJJNh+rpsnZdCe2uEj/1UC0Ak6lT+Ap432
aiEzWzVkDsnt9NQKKceqPsrkqntHzDFz7CDkKeTkm8c/IL1tdDSDpggc2FZM0q2h
q5wEQ8elGFCWXvpheumBtHVIY4mr7oueVCm5Ursi0zHyhxYQkqpldV1S3sEslZAz
adjLwUgfHfEVplbf5WGh6ugAv3K1qy31DxbXHkxOQ1WLhohR6/YBWh8tMb5HkbGN
pLXxBu+m4yulLLiwXnE9uKxHVoTVn9XtjMzX63WtHJr8j6WA85/Voxdb4t8GZqgT
Sj2xGgf3SyVefahrVl8dv0NyELAWEef1eOw96LonVppJ6qNQL1b0x7BImIPmdTbP
MYGvCaoV7i2ymJoypRaqdvUhJMpW1TVhv6d2Vc3roskZ83rh7T29HECYZCSKvRtH
ktmZD7+dYnJS5htoUzp/kvdYIYbrHRVvuQo+8Uboqt7nM4IQie4ugHRudmOBhxql
YmCJlyhNay4Iamso1FQLz2B9JyfgXZpjwUvFZTlfIF6ByLjUpHOEtSvA30Hw7ri3
xjWRmcIhEkcbjUvbTSNPDKFnwyxRs4zxEWGfAtOaQtDd+ONWUJVB1nMbGgFWLfbz
TmBGWSYGblz1kkiWfrkGYajk0SUJTrwtIF41Cm5pnMhdQn6RL/Q7cF1vg6flWWJw
aN5WPlmR1aUn2c/ckSe/FvnpnZ3syBZvGe617EM2dE3KaU/SwVDGjRXIqDPe6kry
IygNBs3FnvjxTwWnT26Vxis7z51iAaSkUIJIGg+asGVcOoEuUas+rIHPVn9tIWS4
SB2gzfrS2EjJMwkKdKZHxeNjaVizuXICGjQoHylRwOBmCa7MfLl2jacUPECNvuIf
Bye87BddHPdg8j3e38In0W0Zy50KEXCOunKf2q59DPnIHytPRyWa5j2wwMh0IqDy
ZfBEOjowqg/t8au/baFQsp6qENQhH5NYhu+kam4eeCEYxfNirDJy5Etp8SR2Oez+
vQ+EtHIMvDXUyScdrp8y+DtgDENkWlzj5Jz0MQNPe+SynDd4foDY3nLrMED46Xyh
FJaRlTiJIIlVJmBfsTQ2S7+QNPH3/8zUcJqZfixGwOsHLc5zTej7RKOZPQpQeMnN
FnmPaKmrSakM+cV0BwxS3/zlGT3f+5kIDNN6ifRkyz/VuDJVOe3+8hn3KnU2xfJt
eJD2Z+lu+LdD1H22AERa2soEuREGWBSzOWDXJIVr8Fi/Fb5L4hLKfXJ8t+06O6/H
DokBEeUrEEwJj+MHsf8266OY6L8D2G96BkNBOEaAcQfTlPiuJDyjIEJgGW4Rt4NM
SIYmP+j8vdQEXCK/sAeV2kIBGNPXh2VujoHPDL5Dxne0zGynkpfbRHqD28cZzXY5
8wCEKDxKqrKdBzbZNCvpZYQ/Rv1k06gtKO6mAixi2WG3MpJoN8bKkubjIHfdLjF8
eQ9P1O+ETYqLIcAsivTR67e66TLDGFPLP0DWnZrGVuMCN61nSsi3aH44+plsyT8F
uE12P8MRGUGHbGz2CATzHctrtouaDgL9WnFPQFZ9/Hjnd+Ocvo/q04mkVKr+UxjB
w+4B1RrZ32JHdNeKBAb/WiJZNb6PQzTFKR0PtcrRu6HlUZskqrfpMK2ti2bEah37
iW8H0vlcrrsGeZaRA+FdiO6awnBxp2rfUwq8RCO3/t1/9Hc0AaPcB1nUsEZQgscr
gUZMSleJh2CTU2tRHEzc3vYg+pnkzUqxd86HDAW73etAAzCdHQ9W3wpcsx/EdGHm
d0jLZnGd5QkJSlcPawfGua2mrrLxkpUAWYgILt2rcpHbEDnXZlbHGs7PGpEOPbwe
k799RanSXHTeDbIAlxIVhY8UsIhgkOg8TnJrx/nXXQiKnRntuyguHOtyAZSecycH
qj5T593ezt/Aw8cVoZx0EpdQVzYNQTbo7G0yOVRY2C5oHSRJ+QmyK/syrpcFLkVj
8Rszz0NoAWHTQnuxyJAlKoVet7dwyzyewK1Hdiv7Tvgvi96vWx89gptGA3Px1TPv
QRDN9Ykv4So30fn9u2LuzGEyo0lyCP1D5ePzYqiZ5m1nZH8RFfO3TYisLzStFrWq
7hH+NpcUUuNlxOVpikSgBpDXuPLN5ViciG6E61iGpKXDIEjxQqzidu5wXttQ2RqP
85h2x98EG+BCF402frii7JbpbT5ek+kndqa8u1mX9hPwDtTQ2C5oB9oarG4ioIyC
CQxzw60/Ms9bIlvpKWDTzpnVPNlSiIv90FWYK5H5vEEGEUX7DfM32PhV0hKGNcrS
UP5j2a7UdNq4emFIsSvhFEKQXEMtna7rKyaSah6HN5OEX8qXcFbnBi31SFwtuVyX
+RvB0nvsezWOuzBbqVpGjQKKbQlrR7vksiEHM0PtfbWyKMFbGG+HEKm82z6FImeW
PEFETY/coWEbvRRBEhW6zOzoAyo2u4iRukUFOBdKynp9n3iwDsGA5DoEUI6Pvccb
wJoIQ0qqz6iTQ9TacT/+K0txF6SqT+AEZQgszzN7/pZ380k4geK2dKpPFOAIu9R+
GHDhQfOH/Yl4ib5V1CxR3e2lxjsWmQ8ZvClYBxr6mjBDFL233OD/WrIZF5YnFL6V
GuhzaH4ZPn9Bd7/U/n1x6HIYYarGsHZGK8JaL/0XHgcsofZelULbn1hPaX+3Hg38
AsIe5NIz0li91k5Z1RvErXCMBzEFlVqBPYwp08I3D54jPELVOuwqfecnQMw5y54t
2zFLGnzqyud4gTBjXCZBAkAaZ/tBZCHL4abK+03EPegvMDwcfJUNhWiLFJXCpnQd
b3RDml3VyaDLrX19dbATGUrq6oCYHv3aE7C1mz6bpxeaDZTDJ1/dhBh6pz/Ch7iz
J2ker/tmgAOruMDD0Skg2uQ9/VIccAJbgiyzZJvkVrPmXnzOVlNuPP6Ea8HJgcAK
sqzNTuxNuU868Px4rhIZofuiqfS8ysjKKlWqXPJohJ1C8QwPy0uHvUBip2wCEbLv
WGCnoF6kRIjK61IICzGoXp0BM4hnPkynly3K2+HiM8FRN/S5WqhpjoGXbh2oZ8Pq
zCDdUnGo4P/jzQtL/u5eZjzI0jLZceU0g8Auyecn1zYvEWucfsNM/V4+yif1m3ZJ
rQomjmpzQTMlUHcX4ZGfWnD0nq2SZpPJDGL7ePLdhoOpx6NrTmygwWcwalaJ9BeM
rY4NddQxi/kWo2ophXqNvvASPJveUhheivFIAk/4cnzCXTImk7Qplz+TUUmdIY61
r4qyWew1/3XQalDKogoV1Cngf16xwSbKIgUFHQrZ1GLAFrcDbXaxd/8G6kC8GZyo
MozsfqqXot9X/XlQykrSfDa8Jfk8EsCwBO6gcEo6xEV27WtN8lUX9q6SiLMfnsEV
Xtnu5gjGxyXup7yuIKnWOAojGIMsibL12pSbNOIaOMq6LDQUwKrwB83oDUSL9eB7
/FK2sW4KSsA0tN7uh8GVSmbFadpE/X84vrdmKVeRl7HfeADIQYlNTauXjR527kD2
wA//DUqRmOC0SGTEpO3xcGaJk83UF0nSDMimSyNKuOq+uwTIEInw0Ohx6z3uZ3D0
gT+6DPEIaKNDKDKict5Vs3ycwKBmjYm4qcSZfTicEQ110HaTpob7JMCkOR2OqpNp
Ucq7XTtAL1QQiXuAGgnIegPx5wVi5llaOA+1XB4Krqbq6w46fuNp7z3aeNSrE/JU
pb16xIeTmkhhpr0ga2ULhOEbqABKzgNpqJ3IMeJlg62rO79tXlpQw4B3461ETro/
eWhQVBsSg1Svo8dPCBxGWDfN64Bn8M7nFH5JPyDfz9NrP5R/DJ+78dG2nnFnixsH
d8+hPm1LIMkx3pO4655R8wzagHcfW0ea4+VT1GKQ4AUo4CnNJGQD27vtxy+P7Q3o
VKc43VDJbNUN4E1HSEjUfRTTi6aTGsj9CWPDLQcT4poH2O09FdANctTMWkml75rv
Ygf7WnonGcF+uQZNvfpaOf5/Z+BibMccyuf3Q4N0GWiK7GXMuzFYAIsvVkmgRYx6
v1sqNalVIcPWgPGBsUQV86Pw98jEjprXXpz5slh8K0fHTlk+sHdE5SwMrhzSsZSL
qQuVxLjmC2bVC0VxH2SGgmb7a0QNNtFlXCFC53RkwW1W+x37ve1j88oPJvx6Pkw8
+HN/ubu7zKrIQ9ElX/Q176KruboONgoFSGzU9o4z9ncO3ivq3OTkd09xRTccjWB5
9FppUsDxWiZGo9XXNpKvCMx3JobAVHak+a36JVdpFnAqW6oDA/e93pyZoPPHKw9O
uFm8etf3b1Sm5hi2jADNt4evhMqVOtxJgcp8BjqKZlaHA0CaKNr3ijToANr4BVM8
NL24sylNeArdFAyUuORUqGKTfR/IGrxR4dbYUPN9UE/M32I0D49NbwxtQ3K8h2Jl
MoFnFo2lDKLl3Dxamj85jIa6nXG/pvZQzbf2291cIxWRmeI+0u+qS1XcwCHUl0HF
Vq3ZpROGPieOXak4qySo2kOw9sYIYNLTykCObVGiwWS9AzZStXup957CTuXWUuFd
IENTSENtrfOCifDwWPY5Vmp4JhyiLaEeLvkrL8OcQropCIyXIUYne26L60YIz+XH
TMk9j7BhM/WAOd8xkfA/LjSReP3o/mP3fNMzuPiHPWEiVs6RUKALIuBqOjhXs0/o
M/UyKO4AvMnnQ3jQAXnNY7k56YikMRvk4TBsAnLoOTSQkyNN6FgZvSblhib3TY5Y
DmjltJM6o6w4qCVM8Qic053NmnDUAdZqwFHoCHX3n6efH1XT1kucspx5hAgJFVL0
+WTY97TWTPPb24R+jORt3Nne9NBfmaZvxlZsLiE3q4PEPD5/Ok3fNuE3PKaoz6XO
e2hEftaSnooqjtKNe5FoupOuJ64+vLKcoRb03T651ONNgowV/mBxetS0ImkjI2WW
ZNX4c/aNQ3UjfiI27IpjuakCvSsu2vvYJwK39aLHIpMg2dHubGgymO2INyK5c0np
NDjy0ySOzGqx0WdcH35qRhQhrcIPewErshDWBCbzElreKAmGj9h/0jV7qBJbRNNf
s95E6jiXgmK3zQ/dNi7dqJiAUxfYUXEM66qhw6ouAfWfCxoGwODiwlyOR9b0sMJm
StXaLZ5+rd2dRortgOUAtd6bGZZXif+Rp2qKa3Mo5m+lgWoI2B+NVvvQyIRCs6iO
ivgU94Acu2s/EQ3bjKD5c0Fk3ghSFZWcAYR9iyrstBXJso4scXELjh9WYsTWwd5b
eNbYAbfmozQTGokMOZzY/wamHmZw/tC+9S5MCmkKM+3Tux+1ahf6bZI+vHGW7M8r
tdMVg0MUhUpWWB1N1B+BLKVWEav1nLt2icK6BZcbgtpmjuM7l5Kuk5/cliKQ802v
e4xW8pE8pFA61MLv0O1jx8gqTIfpBZgeAIhTIvNqr3p7ozFGCILI4yV6o/8PO0y9
FB/qJGBjnB5pc5UfNm26biOajQuGKiPU6Obbk/eLRyW1HVjf5yMpkpjry8prbVC4
LSY6zmWlUr2mrxOZ02oVo8AqzGZJipVJaIUml5knnMPAVTrwHvvaEJDCRNKOImP2
hQ2XaX5J0r+k8A4M8AdheS1KLKG3zmzSkOOwlfEKamLX77usXVwggEFl5RRLTfoB
uJGZ9ZoWx9oFQo6YRG/27BeZ6jLa3gKtEZx+bdZVrd5HFNMpW+yHsD3MlddojgBQ
qYubUFgq5Xdy9CKysWerzoDk8hwziiYFhhPqt1wENhhMDVacQihuCiqSurlZeiIB
5QV/QgGMP/eQxZHNaNFXu54IkEKisSi9o/H9o3MwsGBD/TBScgNna+86s1kJDz6e
s8XuvXDZsA6oKHK2uDKJrJdSB274G9nWAnrrEbIYC5UPm2n5c4OMQ5+Qz+Of2pDr
Zr22ROsdNpySQcdtir27EGqFLKYofF4xs6OJ3cy8G7fa0nqYDbLhMcTiW3npEMYY
jOCixdI+Vq4VBAtHYjGUvQCUHVqmOtIDg5ioAMLQ8ukxjq2NVuyZJR+ntQ+CWIOY
34HjGu22rckhhVhUlWRV/zdh28QMiER6E/v0RixPPQaFDMQ/bSzpuw2zTJDn5d0P
TRmT3xZuUUbxT4O7ZCfIBvlK7HEmPgcXw+IDoFjTrDygp3JNcnBdiLs/Nwx4rg3Y
mRu0wTdoAy5wk/cD9kSuTzeCb2fRwnwvCwE3PsXk/rji4eHjd1HfP5t1TSfNP5y5
hfbOEh9Z00aJjnRqv82Ef6fEkH8B8ODwvofNkSw64vGxEJyzqY131ON4hnPtY41Q
PQUsJf70bQY0K5RA7IdFEvVqGUwJAPDqAeKWu6RmEGasIh2KVTtdlxRHiB6IKbYW
xR1ONXU4IF1TecipHKZ1F3bZJZlLCGFED3xb8S0ZY11o4HnmbuYUcaDyvS/OySuJ
X4VzH2WjdjNVsjjfF2rRmMmlwqhJ1PQa7a4PLoz4SBOnqnwb8hbE15DwDzAIz2WR
Ds+a0qu+3gfBkXE+5lY0uHcTwZTI8aDVWeWXe5phzqTsTchzUPms13cnf03+Sh7S
6g8+FFBQJG0HeLdeWe3Zj9OFun72T4ANXe78GaH6y5pHOfGg3waHoEgtlqJr2uhI
JXpolZAuUPEi0pSTtuo/wWdHIPFt+w4oDCZQTnkAwABgTIXIlCkTpzbsC4+JrcOz
G5YRqwtnHgHoTSgY909H9hbaVLCww/e1JNV45rmKF+cgxUvcoScumKJ6hVR7KmAy
46xLFtED4c8uh/G9wJSAi5LYjNOz81ZEVZprQx0igxICQhlm2XVtgjkW0Dex3kR7
opXl2CZU4pgXveggmfpZoQNkrZ92GtDDpzcc4KOt8KcQiwYS/s/4qT8QMbVJ6HgO
iEOXab5bi1mIwUywfz3SXxCPreUS+KJ0VAsDmScTVE/lpyalvMiJaPp8DjQPhqiy
zxjtPlT8pRmFy4Lb6l5OCKdSh3juyxfwnczVMl9bSeefqBrvI/QTQ2Vq86cKHqV/
NY/xbNRQLOPN/wdumbqHJzv/xitGJdFgFiVKdMzWntx1rlfp+Lnn5qi/9Zz2Adii
qK6Bt7DBSRTeSsWxsAOtNFAmn1iwfr0kRYOx97uFW0KRqG83FnJFTjOJfXc0lmNr
9OUim7j99bq/+cbxTo2idE+Z2Ju/NjH8Zu4Q4zzUS4gKpak6NIJ0E3c+t8ipP5v9
XM60hXSssPkLkUlafxwv2OM5b+C6RjsrNpCPZOjbtVjn9xX1CfIMASRSCdxQwKnU
xJ0fBX0RY8mqkDzRxlfvWp5rGOpE7ZJR3ii7AqLirDHwpE2qRJdzXMSX0ZR0V4ci
obwl3w/CWN53QKt16+ZCyIVI8p0o3szpWRAEzUhI6Yh7ad+VGKJybH/9kYIpTKcl
r2fIXhrPRXBx8E0Q+76CJ2k6OrKmj5ueqUwDuVPctiWkJ8QD4R0prN1PIM3C4oPT
ADy6oD+xo9JsOQMqXJqd6xPmNDTC2VqvygXHiV68Zc+gIzWPyEVyy5ZdEcL8vxld
oSpfAvTxyTajHE+QoAEOWoWmEzSaj1Dn5J/3dPyKqzpoqeghmvTfn4Fgn1fYv7ZN
KzOP+y0axCcQEctDF2m1A2JUHHGMyFO31JJjVbnNbWn7V18Aqb0cRFfRpQB7nZ09
hX3xlLs+MpsPfgVDgiLlMZPaI4unDeQlXZa24lFpMMXIWyVf1vQmYoo7ZAO79ac8
UGk0FmexzbhRqy5Xpd4oybdCGXJ3HURtWOT7o2fNfCDOpOh3g84WaTn5hsIkstpi
uR5jfixYJpHTWZCobAEu/hQm4t6j72GrNSe3uwkcVineWypiVANbi0gJdy22PSUQ
OvhDPMA2Pi/JmqsKc0Wa5vPsoR5PjvHkju9ghC8SXNHaUgrPL4JeMpKHnquZ69ik
lH+/5red680Zfxw8NLwjyJt0pz4fvSp3qYEBv8A6iZLn8JLtTNLVWvlhfLZHzpzZ
qzXY+9Ty0b9pJYnKvJGl/8DZeZWshTqC+i7W9GhESBiq9jo9zULtuYvDDTCilBPN
cfEwn8HHeIPZqj0JA14kVffHEAlxKDK5y/Sk7qlfKIJPgTt0uFjdoNagqkIT4N+S
2Gqikk59a/LiboqagO2H4PuoPRuaHnWr7TEe6+8+Axz1cO5ajHMJSc5iNtxQz9eY
7L7LYMTqRErPhEqELSAA7VVr2+xuleeO64tcB0nxNrivvnF/d/OnE0N8QIKTGAcx
Wcs/ILg8PcZieesuAVoAzkSCj6jxRhQUjS52Im5Q6AT45yhaP6tHRKW0n2mP0L8L
FHrKSIhrDQwgLAThnLzCqz8VI4cxw4+VwNYORxrWMPXOzNQkkpgxUkfAOdAjre+Z
YWkgHpOhuzY/zbyI9RhGUwmy59yBGbHh9GMc0a/vP6CGrQ4bvRS0NWDqWOMvXzlI
fwz6R4ptNJY8Y5Nu8qC0RuS2N0/HININr878B5uVCiiZYCEoVUwusebMpPN3G/7a
SaC4sVvpT+SLZhGQMqXHnM669w5yGmlHwEJ4OP4kACRc7Dgc2m/Z0CqnXk63zRKC
ZkmWF2X4VI9R/e0bWSf8F67jLn5FC9Lm7Un5iY0v0mSilIvwFkeSFVbr70cz05uy
44J11ukER88ZoTclZJCAscCGNxW5QoW5k+rmHgqxFu2Np1ALAMoeBDRg14wOfA4M
1U9ShyAvwz1g9OGWzBWb014hIvPOCuvcMNMRGelywAwIwy7+eR061t2Uu1wCG4MY
DpZO6guQqNyBFmlGuzNusrBWx6artkTDZP4LIsq0o0JybXvudUvyUWhCQEINoJeH
5bWTp1dL8hutorEQpSgxsZaeKxD6xUSGD9LNWd8vRnw6/IR7/VQLVa1njlG8pnUZ
CwZphWaC2V+NQiwGYuk0E91wAIKges0kSHiCG6uX01MfeXCGUs2Ccdu74cZcPbK0
LJzSeM+pN5ZamjXCvnErZEmmswz7DsoHuaZps0FFD9nuPTc7vCAgXPCYOesnZYmF
JJ50h8yazuSEoDeql/AL8liwBiQsb/9RJcPU+0mugnwe/lBisCBJuT7jyJucgtrl
e+d3HuaVnb42LrZAoM0d48oeEX9+37K1bWCSsdsxYJJW9ItSFUEqN9zeyTblTZI1
pvrV5WMttWu9FtV9KQS2jfPNdKDx5qGrnnDRsUdn8+UQRChK4IUiSfDkraz5hsLs
PIMTkC9JM52uf1gRuI91BUfDojDnSAZAuh5l0W3CUDHBMxIKpObfN+S18b7czH42
WiDVvKv78sBfZmebfzklTWwYpuCS/e1nAP7CdNWEfrKSDUsMqswqBWipkd/VgGj5
yYsAu3AWDjfzAbDokHWxgOucAGkjS5PHZVcUgRLvtKQ9OrD7lzzWIcTiWbNjRKQE
bz29VlYzkF+tUHab2IccvR+QquxVdKvYHQSWVQURZtjyKDxCCeh4qvugNIVfQsEg
KhtRou89Df54sR6ObE+Jo264zyGiKWZiZF79+gC0k61Dw+dr824Yk38ILAcUST7y
h2RTGmMuIe/a6uCEUqjLUxzV70tv1cvr+nTeAo5889bVQGPNoOI7pOl3o0fZrTlY
/63cxg7GYKXV5SEMxZIydhbKGw74ES+4JYdHHtsxX8rAbrMd0h98AkaM3cX/j/A0
RBxzB6HFVmGFsHv4TMlg9TcoauwuA9hxgiVQ5pvoloDRvIXdfTQrM5+mM3X3OR4l
Asd7T7ZwxFerEz5MRzcNyKU+PHwZdQzZGE+P4tCHTsj19GqFEFC0O1whkRwE+F+w
R0M6ywEUDv+UuGnEu7s+yPx7/s78+pYEdrbLuTAlrqxqZqesmnxBYHMfRoGFgsGg
rdXKK/nGkepIWwcngQXDN0bgyaZavFFf/kf7iEtWJmI5ITdAJqg1/ihFubl+DkiS
XQKP+y0tVEnxcbdKk8xrYKY3801v9aXoqsR69eP2jKoKLFCv7hyTsktUY4Ax7X8V
Xu5n0LQcBZoIbdIeiWqxkKvg6OsC8GoMoKYGmPxWDeQk4BqNkylLT0DSkq6Jk/3x
F8vMdPNFBZMs8oTDxNZjqm9QVtZs1tCVveKfb/zJuEdNNyGr5KovUMhCfu6gkxo/
WTPIqgPEf+Fhwk8lWPrvZX7G/ppmOD0AeU//pubNeIn3YgvfZNOUianX0XLp3K3D
RUpaCddbeYdfhjid6BtH9agb7qBgFX7qUuXgV+LIKBdgYKLYO1osS1dn3Vl9thHY
YV0yMr/CMKHibyIOHl7R1ZDhQJiYU/gQIO7GfiFesI82Z11n2NYLj94J4CPCt6xH
SbzkeocpRJdVCoIetm7MRKQKB6tjRCYYlBP7Kji5dpGPfB0O+zTHaomfIDRi2epi
kHkv4yXAT6ex/YBHJCcLORFm5kuPazUEKQKW2kqC3HkN/DrY7Q+Vj/ooQ7Agp2FV
r1RKxVuld9vWhnrDMhhJSDEJxr3+XaN0tYWOihGrp3IIudT+hbZgPfhcdOd1IfMT
SzvxnrLKMo+OjoE4c2Dmo1gaL03fyiVf3mOrFvZNL2rQOsUvpY7GfwH2r8xCHjfu
UTfRIudfAquf+n9JK4Co0xsHnI2/8lsTcaPbMvZypL5R7/Hyjh+mj+fLdeBfHHc4
Kn5xsMymhKnFajeEB41unSt5KURjsYzhkJZqaRXNRm7Kj+rjaprF4WJpnDrmQ01K
/3lIm0PQL+oCta9q5XrNQVnhVJN0T4qRDrJdUHoBbsONHi+W3hIWX/NXLFD5ALpl
dBQxg2o3Oa1SVWS7XnLCSIiDhU+umTsqsCtQh9b/nUma7BERXxEDzg34ht9uLvdQ
GQc6U4tFFtWt9aE6F1lby+rc/NGaN9e9+eAEhOvBA+fMCX2XzEG/4BAVNLJ4g8T9
3mXXsWdU3CWbEClm/+jO2/bv6AcfVwhvj5rnZaDD1TWPSVx8nd2rpgP8iLYS/6v/
tRkwjJblyUPyP3MfcMFGJQQI1s3Lnm6Y/Wfl3BOlJHZ10fZNaSrSh6G0U+B7z4h3
kJP4mfVYPELrTcTxo64Dbw0yAYL1L+yeSK1M/6yYGObwLU2L86fz/b3nS3xrG5wE
ZLQn3K1/adhc9yl0xyz3ZxxCQ9ANvxk9PM7yyxYLAK+dJtDzrvQKpdp6fabaRBIW
zTuNk4CbkPgs0bMTB2Vc4eA56SCLltizxdM+mwD3rj+X4EBXKJ1FpMOKj+0qjncF
accMltGmda712zhqZ5DS1VUVGacI5k1XCRBIXMvJngQqDEymxTXB7wxZHfp8l9gK
MqmggsTCTAPUIzHzlePk0+R0Sl/S8x5RVfkW+G1hppJXnh1ou3xL5M+MiKi014oi
rnSpd63kfdPwULwd8k6wbTbd3k9NT1vmK02uOeTGMsTqe+scqiDYzfmdTOsjyxgJ
rq2B9hS2YAgBRaVLqNcYULsn6cPyskPk0+h2lJ2FEaJTRRwycxwBPIPqW4wlpyLE
eHrinjQ/7pLaGMKgumhST8g8c+N+SwXDkR48GWw1lgQ9bpcKigpgcZ0KJJWUC026
rlANW09NYsXE9OQo5mXo6dIzIQ3SmqzvpdIZYPAqEaRnvv2BoVm1tSVJKopUs2/r
wXR5kfx9nKIFe23OwqWv+buu9CZZODrDhraPUPgo5IcS8ixIL7tRKee9fsOf3rKY
n6A6M/DpogMjArIm9rvZuNqIhBfkbKQYmS+NQN39vlq1FtqmuKm6FeKCq13EMooc
K+iRFroI8f3HaSG/8AYCKnfDN5vubgvRtLYg9IE10lahO3oHjXPjZgAwPIgBMD8n
q+D2lHdH0k+9q7tKelqJkkGg9lhGoiZfJoLR7+Kg9NY3YERXZEev3iwurJmLpjfc
2imafxndV2jIU7coB79YJaqHwz+6nzl0DqiRExwtiNCFFlVEb0ElfAqUIwyw2Hzz
ITLzohlUk12S2z823PPdwTQYqzIgYd1jdbYUldffqoiZju+9menxjjotc6lD51lg
+r+0KlveaxMzWqFIkZC8v8+PMdej0/Rpq0BF8ymo9KMqDmqZ5OKDpA2mJmiDX4zC
pAhQcD0rg+YQ6CI/qfA2V92sric0yVB1oNXX/NBXnelAB3K/CTxFQHwAtscLWv/s
upCxRBiwX6Bfd9CosgmpRQeni/vJjiBnSnP2zrgTeoBJnNPjDWdAKtZtY59EakUE
TbVqj02sICJ2lfo9hhTB7zivxNczJHEL86196IlbxAl6eW/LiQqT+BFkhAZVhZ6S
kkUFPi/Do4+gldbVRPUqIhjOsOfqekjMKc2uOP3GtWxNnmeMfUHi/4K5Dqbszu3I
rXwrc0IAAEgTlULI1QHMkaNdUfwp0W7iojPHtZ2wB/30eCSmlLGbsIXEPYt2VcR8
RHPY4XGSJ1NAktjs0Xd02fi0rFD3wztOXJPrx1GwJdjpVunHUxnLRKhQb2A2bvab
6zapuNj+TJTDb3a3Cr61N0LEnAvMJAFibAoBG4mVAe/61edcq8+zk4CTks3K1/py
0Fmcvm6EN2xF+D0XnR0BWuYAxNC3TvR38AbwOr3S2Mo5zIbqQVRV3Ris6vlNZ35o
2mteqK2ci7e/BI/BSquPdrAIasN5BjZg24VBcmZ6SfqiP+ho08RXZJh8jRNBVRz5
CWBVmlJVzDlHTdxxOE4cLioGUu5TLnv+8m4lU1XeR37dHSojlXammbWdCxyVBU7Z
G+XAILIRU5nOVcP0w75S5SXKaBFVbq3SRVxmg4kn+/odO1AfshDu41vE+DpoO0+5
`pragma protect end_protected

`endif // `ifndef _VF_AXI_SLV_RESP_CB_SV_


