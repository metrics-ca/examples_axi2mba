//----------------------------------------------------------------------
/**
 * @file vf_perf.sv
 * @brief Defines VF performance data class.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_PERF_SV_
`define _VF_PERF_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
IVgEf5buKy8T9UkdyxxNVg2hhnxJo3Cftwz+AV1KGFccxIq5y1AmwdhGA7NHKjGA
rJ1G7JWjW7prj0eMD+IZFDa3AQ4Prz6PUHCfoXyE7X1aeQ6GWzmEjxoERLrK8fJC
sAkcedNpnvvI5g+l2qAAhuG/YZBhvyjnMVE/3zWlWHf7v7e8t+564ioLEuRsUEj7
vUVUF4s4+yjCXCZi8QooW/Sx80LjAW6Hg/930Rixj8s8sfqWKOKKFGZbyC57YDR2
UADD4zfmYKlQKhGJeVBuACkkC/aospyjdsYWuBYag891ymuKWEf7N6qfs4yC/R51
dnczF5rANNwmRgcFfeSkBQ==
`pragma protect data_block
whlRItwnCrALuugf4mKupEavKSBPvKk8vguyy6EiiBY+n/0FR0/bIlKZ4Vgc5NTU
6USg0bIcuy0E7F0yZE5t288g3PlKM9sZoUg1rKQ2+TwZmR0rvTgnoWu6DuXj3lI9
dihB4JgkuFdABbOeFlU6jQZtObUmTm+tsC3wuCcqB18L1fA5m3jpD5vn6zS+ZVMl
b9xyQZio5K3n8oxbhlb8kqyZV2WTO8we75ydAcdd7dnK5rfcDceqMks8Btkqvmvn
7eSQehw8UEpyB8PVEtK8rHMBXyRPsN2FW4Vp9h5Cs2A2iGcpQUELgB3xQiQu6Pqd
h4KUBBZFNCVWZOw85Q6h6px97rsZ0wW6a3LRC3yBdbDabHOfarbgPEfySxGlprFM
PD10UpD59OCT/6hha5NG53H8zVKet6pCwYiRSdBoM0tl8cbm9VmPYN1mvyYhJHiv
acgOv86KCk0+P0hRFrbH4fxXpcMTcBYy70PSZ2UmWC+0EYgfEeDcKlPgaCGCFRuB
Azmu12/kIs61R1rTaK56yfN94dUujvk/FQWfUJe1acsWhbJNbJNb5Mfn74xLRzvb
1zUju2gXqgGefL/4eLFITU7f/SAOEDxdeHvAoQIO0aDafDOx9opWvEvJzt1Fa7UO
vxABJcppWIlrP1WD3AFMmfIfn5ySiSJKGgf6wZEHTBOBd8+iTtBeXfpmLVNdz6H6
OIPscK7KAu4kD6Hlh5qA10/Eob+kaF9QTBF4pWmyyO9SGob1W9bDhRmXMINlsesp
S3rhTyOtrpronwIaYD6tGr3iaqT38xu/bFaTRLh0oNFaa8OxirAlj9B8PT042ard
CAJ1JeZg9cxZUOLl9YOg2aqWAS+6RjHpl49lq12M+6enKQ9UxwTNTmmluHkrgmA5
Jz5G4YC7IynBEk3/k82hOWEW0rnp08G8cjHdatp3Zn8hVnqVu8KEPmulB0ssBIHP
qG3zMk7E6ghIbx3UiHBnY6lMBBipQoAEWqeND/+81xPp/xIPCpLmTyQgkVvch2Z5
D3cs0QRLssuYZG1USpyXu6Vf71TuW8mtd5qVpgiwS6EZysKZwb5M75D0NOXVpoUO
kvA4VKulmVUCsWa+AFxALvtfL5eETY4rK2yJWk+esbICaAS+2INOm1xl5NexfEqO
Cixo8BTS9qRBZHzrslFene3VBZNd6zsv3qkW5hT13WbnahjQMjJGYDGoLomZUQXC
eFzwPIQF2Ud09A8o6qfe/b+PVqA/IuvDMgBM5VhN00MdEuPnNGFiHn1x19ixxvrv
9iGNRl+F7CPAI3efK4dCp6JlOjAk9lJg+OGZzEibFQ3S7b8V4vKCEDqlIRHLa0FN
iJSzmGUYw0euFMZfQWg4ahhxxwAFr4LGxexrlvzbFt5dd/2x12ls6dtjsAerE9rj
PEChnSWHypLNeA1Zu9QxcFJjGHjRoJa+1P0rB1CRkbPNCiKe8e26fKZ02uRFxPaP
hrCqeQ/GqC8I04U/HYZMMhtDzmLb+btFw9dGUwffUNFYD1AdgyivZCXCPm/bki6/
KaUKPTzmyOb2C+Pt8JZyhJSNp+Xa9JiNOZuKd4lQ/074hV0kiezYFMz++S/UHLPc
p4q6nNtYCgiKWHQjLzNqZOAH2JJbfdNGqxyQeKKIqnxrQ3iBVLFTzExJ7YCtKJwE
KBMpQT/1hA0JExjyRubyHeV/zL/rtinOd22zgFufxX5tW2vMft7G0EKNCN+pfKtl
DRGOQSBezj/BtdflknpXtbMA8a+hwKDFL5kzlJr81sK/ocJsJpkjh5VGpq02pqUR
j8VKMhjsR0eIlzJFcB/Eb1eKWd7fmb9z7tzEkVyW0Po7a955BAUvg00J+gNZgXuC
Mzlsfj1KoZVG/dsSaOu7sD1PCF9DdvYxEvvwZsA6rl0jXvn+/nFzJpfEv6n2U02a
KlNq5VHXHLsRZkQy2xN4zGKMkk90OxEEABV6XqqUcjb2beOMTYCOcc7n/TBz+DAE
vxC2rX+oRzftQBxJs+QlP/QC/vUTzVfCcj0k7Py7kim6eYTcf9DNv0eebuDVmvHF
PYJ3qwFl/6FVVYanZchJroEYC+5D7ypioirqQYSGkL50huC13e05/UEZfQs4+lty
vl9Ilr93eqpJYUu90NQ4HjtpML5z/+mH5cmt3b/TAgB3xJw6OT5yJG1zEFrTYsfu
11fMpUhn442GCe/Y2hQJ4a9stpfe29BdQO5NuQfk+R54IkI+4cRvd4oIp8/mN0CO
+97AbIvNKFsW8nRaZfzGRMngD/wNc/NE7quS/Yj0ZgvI3/WOk82jSqAH4nx+MPq/
gYqOBMmmmA6ishO3/ZAA1o/qY2qjao9BNvE38KRNUy+HS4tnmQDXYWLdXOGPijg2
gw5Rfpwk0DhAc8dSNiCohkB1EAaRyHLgI+v7vs2hfKySvqT+9UC2EJRRlMQ658N9
HA5gi5RzsTmDmfKhAyx17BgBUC8zk6qR0GvvGT/fsTu93UEMVGC30a+A+UyiBP6G
evfjSR6eOSyauUrkFFUhFDspWF1a385V8TDtpO9h2uMm4Nr7zuhUTp2UInF7rpuT
q+hWzS8CVLPZwOTXLyKk3LAhVqQ/MtjKidiOY0peGx5fvz0oBVHlFwreXhte29GP
P4MFi+PkICKtNXix8aS/X9HqSGn1NH8/cCkAlU9mCVbIFSl2H+LQff2LSCthDo4V
6oxYuGFBYgiuXa6T7lKCTEISQJwu2QOUyV4uzm5sxFqYmh6EmYxQVeDH+viS454x
iwiVpA1ncXY90ySSqpR0c4KEnQDxBbZxaiVj8uyFuqy0BhRLcjaYQ1Dm2xQFpoEJ
m00g0LyvhzFHTgDVPwUWLLb8/y/WEqp3BdE0BGgI6+JWMBxmhcfuXcHJbEh6YpV3
XrlwcY24VPHloXUepRH6r6Gn9SXg+oiixSyRU+1LNdd9cI+4TayIH0DMhgaI8lZ9
1rEEHRFKIKyKcqvhstFBYnVFjM0cFlF3dI2SaPYKazgpg2WTgcRrqxQ+2VChG32r
d+Sc5iAu1b7E7qiOuOhIIYXdVhsacylqBrw7YxvRLP9piXTbYUzS94/1saKvirDt
FGAiotsbX6El+LS41SSZd+A2hsuaCcFhKKHjtArc+TPGYeVbT7cdUzB5PfOMjWCZ
DOWisQ8KtuT76WDdiVnv2K/vuAbYmQsqhlpqvRucLBo05AhUTdrNCC0Yqj2nXusU
g8WegRfm467TkTuBSAhARb28wE02NS1vtbNsQc9KbU3cyRh48fymXIVAlhT0XoJQ
vfDoNArqqpwPFxFEF9d5wbpsxELGWyq6gNEZkbyeWU016Pjm6bTN3qKWxfDQ9ar1
cv/tzrhcxWtXUFp/StuvdJHp/hNMUbpjUoWfKmzsFyNyOLr2eyXK9Z8xc8wCp2Yj
3jLaSfwE9YBHjdbI8NSJ3+ZYW24TTZRJ5lZHdhtYlBxPzDTDznagTtlKkvGsAGuW
+jposrKrKVhT8MTsrnhuCDEqlMPgsjRKMICoteRbctnUvQ0UsEPW3S9bSAz/OJcV
DaJlUr+HQoTjVcaXbdwYAxyg6KX2/3A5qDaK9iM6VBN24+R59QUeT4oqjO1JbVgO
TS6GvFuE+Jzh4m4CJV4zVywdXc7f0HVUy9sxtgYi/4dXETTYjYR6zEGETH9qqSku
QetJ0A0Z8xM5BcVmX3Rx8QPTwIWRD0UQWGQhppu70tBk4pUt/oVsEPSk8Fyd7yhY
+uLbsZZvTgobiVYvIE0jk4AORzXZf4V4D9DlFzQ+jyAz4jER0GASKXA3ov3Y/Otq
711PFK6iHLkltbmyc0QGV3IfE+f/HJllL25lGjDDtHx+5i65zE12a5mK/uXyZ16j
5OCURpxp3Q5h5xQcP1Zg6FgPyXu7oNkuSVWq4F8tY7WzJ7SMxZwRD82MNAcOHMkT
5Tpcr8vIB0tTZJJDUr9lpZMBPzo/SE40Ep7AKubsyoJSdZQF9sj5vGaKJSbLJfVF
uXCweBn9weKdcYW/oDmUYVNWyuWVrkcGYaOd6xR+o3wQED/ag2+OsccdTHZASheF
UyBR6obsi6T0/g75jjZJvi+YSbedpQGuWcetdBZSFdWRAB7exSRqXH4ghuKm0DDI
fBaUQVF0vD/ZR/ZdNrvxv8RoK+/4hqdOgxkLg+1U29AOwSoY4XIF9gCFNR3JVyVB
O6QwUsGgRY9fcmOajAdiirKU4csr9KflU3mbIfStk0SwEKJGWamdPd+WHfA48gg0
w5+lg+NgehG93jzQn9WVtRMbeSmRHXAM+Lz59N2v4r092i8BFyvng252ydwA4uMd
Vylszqnv0kXXCrH3lwts1HaqR1yn+6iEjJgcdmRaOzgbts++hXBp101Khg+Lwkid
dfttT0IyiBdvm0j+1bhOP7p2K1xpNclX+rJ3bd/8JeQh88zhuWR2QvsUIhaqyp0B
lxh+q0emFnbpQmh1wHiMWEWCsyXqTQL/KtNhTIHWAp5L6FmpVCTOKArzSRykX6b0
YQlK7edbzg2KV/+I6PcOCNRnEIgEI/hWRniCakMXz3EN3UxUxYvZnQBzk7lyrxxZ
GZZ0OfhIYUYeu9x/bA9jxZD9jjqgFxRIAZbaIhsN7cowXegBM6kIi/m6R3TdBfjh
GkqFpcWEUI9M2iqzxFrgIkAMR2JQz2fQOx8Obcc9NJM4TqvXY3BWJPTZlo7xZ6ss
Z0ckQ6QLvE+5QX901SMw8QI+tnGrV0GTcBDLdvCBhPYT3HxCOjTnsIdex/YxFINZ
zP6jrlQY7RzwlWRhZTs4lIvQYgWILVoIDkhn+lajT8DYL0xflCxWnBQtj98WOrH+
3+yl5ZSf8J+yIAUEReyeVvmToSTlN7ZFgdsSdJ5DKwXrUEF0FRrjlUV/dK0m+tjQ
6akEZj7VP6q2cD5EM4dmVWTXa1uM3C4bdhpfCtyzJv/kWmw4rM7rMIfWc3iCq7Ff
AG8lcVWKUxpEjELSzKjPmiii2ooANQBWbHXtY+HiWtlaGf7M8fL94f8XfICr9EGb
vcoYZ/ymwk0lTukF0AqDdwtDxxXedd0ZUl+AAbJGh9+8pI6i3Vq3W5n75RqkeRJb
54MvSYMs4Js/GiSkawXlYGgljfrhgFj+qloYvkGAFRGmD15QzEct89Mkug2LP7Ko
OUDnybGoAgkndHsML1Lq22gDvKK8zMYPXnx44b9LTxjU/PKgy4eC4dMxthcHXfqy
FsVRUl9HQFazFeWvNbn+qWJSMaNkPviseiGWdDuit91KSkDuaYtKC89Mu53hb8pM
ZagDLdXa5uf8AowLMUAU8ysdrsY69xE7rupiToWN3rns8BOysNDFx6tCtbRNGA8D
/e1TWTsPyOIAUu+AmzZukslhSpjiqeRNpQyBDmMsQYPRpmI7sQKD/KpI/owNBZ4/
A6MmWOIrar9nUyWtYhN1z3A1BhYbNvFmtzMqpjJ5fVgrOj7qIFO+lfYHEbxurklX
0khIc18vQaX4i8izaaRzsUlW4Oqa6ZquTOC1BOk9r+SJbKluGFqOubUoJPTH9G14
MUsIiyI9ALeB8395a4Qw1iDN6dbUYQ5gfWy2zd+b2n4Vd/BQsDkaIfSNYkL+BqzT
I9zkpvfy9SOxt3E6iC8EWNOidVBUr6FJfHZ4JFiCXTq9rAYRTIJf1FeZtUztrH6/
j+QQo+2Z4j0lrs34GDiSZpcKidxJNPAq00/b9PyI/1JVV71w9vzqOFfHTZ6ZMwwE
ntsStJg5OfGGWh90299/z7XcNrRTS5s4Y/1JdBxPde0SgKO/I8bZDywAOYSqPcUR
s4lRGkK5RXsUVKgp3aDKviSu6I3c4Y3ShH3hfhUhRntZYmZHqE4j3eH4ThG22qFc
xxUdDctdfEV1UK6WlYhD0QAQ5ONVoMEGNn4357BvP3KjQYqnrzRzoWe7FsI5/YCY
jGLQ8M8xFKOsum6R9G5PKFCDGObQuch5PMhzU10cML7yUNqbI6OH9zBMBQl8D0bb
PBQ06D7Js5R37ELsZsRZRSJZbGwLVyah5v4WTgxpNV/nFERb0XTGq/JMJVTZdqbd
rzxTvERE9qAcIbFlBeFylK2QksGVoRrFb5TlZPTo6EKNOr0uEj62m0Q5QzypTlFN
H5V4rDRpnqqhCIbF2G7jGYUDop2B10Ayhsae56MddYGM7sAS0Fg8YQADZsZZ1Sq4
XO6OkEpuhgVyRmy9NqLdpNLRR2bti8r0tLn/fjky0JtsL6yz7wLSDMPwmwNhTdKy
rTOLIYk+4uXta0oUyaT2QTT8lERCQaJv478NskJ+Y755nrEM1/eaQEjjtSPuaxQc
apQaftAJPWIiSlj4Bd2FXghlAuh5SOwtEYGBFOBgL6uW2ywwreQOjpx5LbKenw6N
mLKgALOOnd8ENzmMAJQ4RxEXEVuOkSuXIZO63X551gMzA66yKxBAPFq9A3nmY8fv
+RAF+37B8hIZZqc3SHGf+M7/j0t+HH4ONDVzTkhN0KwOl3VU3unjZ15YDUbBfMu+
W8bvX+hLiPxn+iYlPYoukyhMqB+GutzRQItTuWEcrOllHkL07Oxj4/Vw8KFqFllc
Sqh+dNV/XVfnxUaiyCT/4T/265SN/HyvhKdLIFOpxqzNLkTWivoUXa0wmaRr2CjF
lv4dMVlOT2DIeOc/jPTzsDF6nNUDmHvkW15SvIP4hU3ueZJb/c4ZhJhS3dYltloS
pRZMh6m7iMZAVbK4HLWEeULjzNJDy7dRAyzq0E+/k7JuRmMR3WiwsNrkOHGp3quZ
lgeS6P8uxgxbhEDbHbuYRtvQu4X9Nt9LyBOr2CgC03fYDCXWLZwDTpHTrAXWXhqm
xn7RGKzOr0wCUG/WtK5GIQYO+sjUDWW8aHalaGfCJfwZEG0tug4nKLbDKb5wX8jd
lPgPqYHKvZYVuPYfRUuaN3SvxbWScsSUbOnUkEdrG5wOwm3iyiY6dcykG5SinUUa
nYMWSUi/qdOstDKvC3uehIwYb4fYu90X6682j4V0oISo9rzBAjAD98QWET8AzxNK
v+OH+tQ+ksfrUeeiStS8knDZFvpzrjAflgtwyo1eKGGG+dUGRfu8cR2GMltoZ5d8
HuGGJKPim3WQHbF9E2843MlcyNduJrRT1nzV7DMvletgZS56bCSVYAqORLbV5uiN
QI/i1ZUB1Zg6dsYTxFOvhRRq7UPj5iJnHBEOJ8O62ZTFjOLgEm0AXQuopWaWT4dk
IJCDiVRGFAnyjDYocRcCW3tRWEC5ryep5VCgp57ZfCTJl8ibxnG0iezRROXlqNOY
f2Od70Vr4/VAfxluioKZNCLS3ofhbVAqinh/pfYYRjnM8BFdnMHBpYGtAFmOpjdi
/QTUa6oHGyrD4flOf8lt6v1X7Sclv6esB98LOdEkuT49nCujEMs3WLFjAGkF2k4K
pMwykKAHwjdhCgx8zTol4G28M/J4Fdgav7UXbs7V2y4tidpwy9+SANHqRbDjOzh/
MLqqO6HBic3ygTGmBgxydd6Bt53AJI9eslfMx/ZfQlCJ+saHPhTTTc6PR00aO/6E
V40qSRbbudLvgho0Ue6MDxH31h5+O7cQ4lRid1tC3PunFsLzyIU0W5/AEthRwCOy
fgykGvk50L2GV4eOz0O0dVciEcNGZznGH0DIEGv6a9SxjceV5dCjyIrXSmMBzFac
wVxrfkAtWVrVdjVG1dVWGT5wulnpe9sQI/aVzER7nYUUYcfU9HrWPLO4r0WCkU4X
hP8edo31RCj5hR+rnA+istccAnzYVOCHL7gNQaIwjM4MCZ2UBI4LDvkHkegUhU6e
EkFpXv1DqYwh8VNMrtlRGOd9pqSfyKNAVqFzp8925qcGvqOtTKUx2SOikAXn0heD
BjunaSOzQ10szcjey6iLvzHSVEd4LRx9Ijc/+pCjuXS2Stycgus+WUXew8S9Ap7B
x2YijOkvkd/doj3erAG9+lmQlxJEuUhoYlICwnU5qAXqiE/pDmN1xMILm0Q2kV1w
xqhKoGe+F6Wf/oBVxwidYXgsE/qvJWkWqgdjsSBfP/G2Z8pU81yls66v/RsBR+eE
BWgoBAMxUmuOKZe7GZ9ApzcQLt9C+djiFolhGfl41b40eJkScscPR8zTt2U/HS1J
13vxgY5e4vDItgUfF2hP2iZTNhxcSXj/fEnof8lDIHwcLDTsY/0kBotUEiw/W0r7
yB6RAvVAMri2Yg9810vCJ/G1fHHtaPLeqhFfZI74/E5hkWBkO99/y5djtbpVC1X5
Nxij8NBTqCOhFPqQWfpkyLbzsDMhGJcjE4Tz4BnQTG1oqfM9ZilTIpxoDhPORhv2
LUA+0fawhvB4DoUPD3UQDdNSqUvmpxe7cS8VmWHKKZaQ8uixE/NdHapayXehdWx2
swfy6LbPg2xfW5eUVNHMKAy+Eol+aVkcadjuFF6GNX/VnbvE5+t5OoEaKi4mEIhK
MDAEWNm8I0IMM3L5SPpjEOnCT8MIdzuuZ3a6I8RbLh65G3MlxRo/PIBhhudP9YrV
oDOLV4CaNHV/OaL8wJkVd0r/ZQzhPlSA89YuN8+sHzzpsAeymSGd+joxUYTBUzLe
6D0Z03GhBqEKNWPCQJ/uFfbTaGVGSYFp088Dn62dugbB0A1373E67dAlJi8qtS0T
xACdEtOpjmWoOv5vBt662dX9KPRKbzKNmuGzGJmtvkggYH5BzdO20e8gnD8mY2Mg
9r/LgN+tCENDODhUetIvlgi9z8Ct+8qFciUBFN8dKqZR2IZWXXJuJuNULCq4tTRP
3VZG2FfPoqWKFhA06+0pSNdft5LcLElEZDCfU3ayslcULNAttOb/foZAndvkerPp
+isWkFt/Chns2nk6MTElqfNDPMcpZO8b1SQEMmMIGlONKX/CANVsas+L8FaWrEZx
AblyjXAY2M1+O175FUE6xEQFDXMoYYscaaORi7hSgvFw2wij7g7FlH8HUDvgIZeG
1cnqHpcK+3L5bK+3hCjSsO/+23jZVDW/c1zNXrORR5/fr+lvWT9qboE3o3UArspY
MY1QFq1fPelaoVzYqUhSgsCKpDJRHF6fu375FhefELK/dkaHnWUJ0WCvYUlSDJGl
mF6RCVKuyW4yYiACwsLN/9J7VgYVvmZzRlaRELvjL4NrOLsc1jt7IXnjVkeabj9k
dFJnfdu2wpQHqH1W0h7mpJKeTtwVHzMEsSPWMSd9iQHRn6quT3eQTcvfQg2GoiY7
p7HrXwtCYf9/ltD5XtVgf7gQtR+aVLzIKjN7cihrr14ccPC5NNbfoeJuU0NNek+q
E1QGWREMiPxP7DLcvejKoR+x7PSlbwYMFG93xhu3m7aykDzV/Uc842u62V3gTUAv
GyEr+fWnLnjATPTSOSntmMKxdm+I+wfXO8jKzG8gTg4qfQo0+Wq2UQdStQgBgjAC
Oq8s6Mq0XJeiRqrq2CRomLJF7FNikG1Yt6c7NrAbHaFXilALfyj9iJ8Y++57WbL4
2rr82Jzv7Ms/LaE0kmMApdqkiEZZDyZnU7VHH4v/ec1EC9aMjaB6wZAAnW4Xwky5
niet8gPZQehAOUKbW9MkViTnmUPRwuduh1FXbADmmm5j7KjI/6GddUCpNZtY6T2q
R2TWTLDdVGfFosFnlY22q5Lr8GjCgmQwz6MUn/ZVfah67JWHezhk/hdG/SM0HHGf
x5MTSoDIcqIg9zxHC61j7ZLL9yxSMUFZqPSU+L1X1SU/RPwVcxS0Hd+erbYVylGv
KjjGVo0Yfpw4YWMWpCuq6Z5AtjWCbRC/NhF3wq2XoqqMwTw5ub9+9bVAiTsih0kh
UYJOXK7lbeoUKRJ+kFnzV2dAjbHf0kPoLyXFxQb+elBXnyBkajwutklTKpDOYacX
lOHIBUMjTMbIoUnbQ151vccreijiUW3hTjaf1ifZklligLOnZ04nTXJEdNwIh9dj
BaYYrotwVHp3HWGBzvE9/bxKz/zgyDGcDx1PXlRVIxhBVQwyplnVYOlPfAwVRrC6
DPkxGGalcx66YEPa6YVD12U+G2N1KZYj+LCGhwwNHnQz0edNtq8Ues51txAEsR/j
JU9RxwX1JvttoLjSv8R7Au1AdN/6Nw2Tw+DAYb2mQwqUqeTr/LxxK73B2cO+LCik
XpyChWqtBHB40kcCclz8uuT1wcgVVBee8QQ9l9/ZbCm5nxXoq35mmDXQ0KRpDbUw
6kjO63v0d1ZytKodpCzKdcxbgiJvWoJ16bXcbdTnKrBWr8qzQI+tA1haqYqGK0IN
rUsE2Vuy8aFLSqsQfxXu7VoueEaPTrbz4KwxbEES7uj3Cp8xtOakFRXQnTzHVH0y
6wYKAL7gp0bSyicEvosGknHNAAxLVrVer0e31GONzdhyI60R+z/RjIf41jkflXBe
0kf2fVJOXpCUbZEjASmH7Q==
`pragma protect end_protected

`endif // `ifndef _VF_PERF_SV_


