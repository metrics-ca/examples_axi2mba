//----------------------------------------------------------------------
/**
 * @file vf_xvip_data.sv
 * @brief Defines XVIP wrap data base class.
 *
 * This file contains the following XVIP data related base classes.
 * - XVIP wrap data base class
 */
/*
 * Copyright (C) 2009 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_XVIP_DATA_SV_
`define _VF_XVIP_DATA_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
j2rJIrEMHfTRl14dLRHfQ4VLG+2j/e8/nUCvAfjY8iXqu3MYtMRsKL2Z91bciMRg
tDwcKJXyTpkXrEFEs4F2T6ySnmxLaoSGl+Iw5sIMdY/o5UysaCGt3wZsqMF1Kp+h
pnQTokA6s6gQTlRKKaDxGZaF3a4wGsHCWlwWHtY/XaWHaGoORnhQv6SwUedXUsp/
4ocwoAlXM005LvATaZIpqgyLVNNfCcdlXL932cKUegNodZPJDBm1QODLnJeWwxe+
lGTWQd/LGaqWJQg/T1cTS3VhGFOJT4tcyxCqTvKBgKoyOZ2+xGP8FUG4lRTt320v
MBXmLDD22aBq0FsPIsBr5w==
`pragma protect data_block
Mmn1OBQa9ziKid5OWgJp46gEvU990mw8xBK+EjdSXKUHdeTw7v8zIqn7oZgBraJB
cOQdlgFJKw+asb1b3UQB7fDsORFFDD7+ktoUnWT7/xHPRpkdMXMFt717BiKsKTJW
4mQaCwhnJZ6xLdOrvz0h1GTW/gRg9HtxdImcz9cFgB+GMfNe8H0ZTuVUoJ8uEK4c
fYxoMey30BeDDfFQzv2y+30pTqwW/dtpJvVf/ZPZj1syMITL8VEBp137JPfI94yy
v4hzZVUgYSqVaFSHRlW+dJQnZIO3Rn1bq7AB4JSR6LLt3enjLoO8+rs6f+Hihep7
S7MsvVuqjswfQpvJCMZtgaM9s8YhzBeoJ/SkfluorGuCYEddjKlYJ1+Q3Pi1/bV1
m9rRtSl3d+rMu1IoEokHISDMH20RgQOFc7LPBJ+hP/m5HhqSVKw54zB96yWi1qkm
aF58IYy8MEwGLdC9bcnbIsUIU4t3Chn8M1i3wUzlUO8nD0sdxeqo1BfA87KmPg7q
P37wJK5NY+C+I3QkMyXs1dX9ozDx06UxYshU8jpw7QAThmnEHn0jQy9Ssqgkcy2A
sB3uPRyLb/i+mssfyCp8BkaJDQspk14HDx1cZ+UY3ogryz/D3+DCTADu2xE7nAIc
8Aja5U74EXoHn7TQ7u/Ds3/id4qiQkbnWTNboq0IZYTeRm7wCPHXokFgUuo6YZmG
IH7zD3ChDQlekyYbuDj/lebvl+jPotT6/BHomfKGPxvOnsCeWaji+bSKhb3DgpME
hGq39qd/kEHKbkuRq67HhutiWjfzdxGvy2w2YLBJheM6HjeQbZXf4Zz2GqRNPSx8
H5rF/WMPdwHYr6ZuFCIcL4rnOurGTa018UbCHSZJ1XkrD+BZ3Pf1FzjT1dsZdCpB
D2UeE28tfH45GMbrbNW376f1ox6p6WbpxqizJ0YGDpBHaV/zYjKWXKId1BCu95QH
31oA+EqzkQlOy3mEC3+v1Rc5qucbXGZ2jMshZLBrH5BvV7KBKB04+6lGhqg/pffh
21BW3NAUSQsNjlw4BJ8JoQe0tBhu4cIENcXHeHQ3w/U7USllEoVdx5xK89yiwNPw
5nlNZPFA+LY0ox4qXZwEbn6a9owYKjyKqjW0jwcsqWoNGyuudwQzeeko1uAc1O20
U6Tu8LSAW+DteCzFSJAxrrFgt3l/g+5gSxCXkwga2stAmH9mj4FJ56L3EDrVog70
hqHweMRD3BV8mbjaqkbGu6k7Bptln4vAun93Lwh28Pl1ESinpHVj+Iee3DDCcUJu
YsqcljK1+ACyx1XnnQnYi5fzJQ/BBFXQlCTAuHIsx6mc8TfhcKEXsvD43H5sdC1F
qPXu0KMVqR+X1TdbfvDcF0t7mSwCSWKLGD+z256jlQZMYYjmH6eLXxXR01p/M3Y3
3eSCRLKQ5iqXPhYgyASwrOi19zYy2nrWXiC+o5L0xNpUDiI0x2QG59oR7OYrJmk0
xqhwQJG7+bPCZRTtXxAYb98UAvUobUssmwUasH/95CSlYAZ6jw1LiGEBWf8x+rTr
e5Pi9GRy6GO+vUNPuXBnhw0NtNGcY/z7xFDXUepKqCZgEthMgF2M+YoNWCmegaby
Ule8R+pgzsmWQT9WkDtU/z6Oe1DtWlnbBOVq3y4+kK90djLhfSDcHTUi6KTqym/j
TJRcNJ179xj+Ey85NWQDVJwFCY6Hg1t3U93B9B24NI3ZSOKsQzr9d1+6EKJO6Zyu
lr5dib/Lxaql5dBYXxt/Kpki0IvsXpQQywX39qUozTBwup4q5DRHoUTvBDHtO+ob
KcaHxAjMD99Z94wFLhvElY+KqClltrCQE/PV7DNMFJltv7WLlmAZew+/izCOtapH
3s5itSoPLheaRoQcf2hJ8Ax1w/aHTVKEVhm8cKFtOy8UYuUbB17kVP1x/HJvzF19
doPVmD1P0hOUs/MvEixhhNpiVx4LCuRoixbubuo/K0N7cQnegUJjWUw2Wiljhcj1
ls3wALjX3NCCLBcoZvK9PK+mieY6qTu7+bvvMuOGlSO3Ml1N6QYN6lcnzVYSE8rG
pYo1eLgbK/o0IQmk2KYX9iOdC3KMVd9iXjEvptcVWldqeun9eJ0bAmYkQH/devG5
EMceaIvQKGMQywkwKsc+0zYuHARXsICZ+m5FSKgv+W1ympiZpwx+Gt/IGf9Rj3pl
y5jz7YaAQPTOrCC/2qTHuuAkf6dE5YFagw1dE0qS+G2I9zUDntW3bJDEddHkaK8x
fQ0mUGS4JsIM5/aXH2ep4wE9H5Zkr2WG/rvI0mG9rcM7ndyjcSTI9uT0Ng88femU
uY0z23+g+po2c7KTNRLMtR1sS8cT+BFcObajgXdncwY/JbRj1S+TYZweBrOPfOv9
zuM8aMquTfkxlhUVcGiBkItMjFgpBfcIYNZmFmXqgyFuNohF3KZmh1L+EBGTaDEg
ZPkD3JO3qL/KGggPpWfxoHjcPKM/ptPQHB/FqbvydtJEkgsa4mCP1H0CjEBJ6odg
DVmapquUOsCxlijmMTfWJzOFhZ002oIouPnS37KFmV9HKu5n6EWF9IgG8S71pP2j
lht/KAPQyMVG0QXgU7ubG2kHxftHB968PVqXoP4UsKAsdNCL0w+HF98Ku4Tf26jP
0fsBAHIk/JZuKPDXYKd47epQuzj0vmBuOnVX9LSFt5fIkkAvVcUKe9hgP9NBpsaP
s8a6CHQeuXejED4JnmNHGsBZTTptdMfo0cC/8hW3Dw7Sc+z8DEVYmnUC92R2YmMe
3Pbu5jyaFyFT5CrSA8fvGv0QY34x53tdbfJ+FFkcrQux7RBIh/70WkzUlV5LR4q4
XzIrZSlsc/Vur8AoHfZm1V8gbwVVBC3FcTAZM47wPEQ4SogJP6wd9B1Yr3HwXA+r
7ukyUjOBSDSbdN9HSRvL6Ql3u+pAZ8GsBf2XbpXkG3iO1+oWI6zqkTGPEFcdtA34
q2rUYfMe4rE7E1Cnh2umMkExmljtueCiArOJd1E5IB2/BjT23kp1rW31VnmCnT6/
FBIC7IzSnMmYRGtUXTRCqVzmF8xMpzRMIllxQgfiy17NiEX9ZidjYi8AqhdP4GKt
otnGGNZ/HAD+wdDzv46Acq84p4UrdXSxi2fiGiqiGkPLRKjqBowXlsMNyo7BT1bk
W4CGcNO3t719xdrSS0O7dk3Z5om/m19yMVYgtc3++9PnmFp8dtuCbEdPZ58PADCZ
C50q2ysLRwJXxhZ7qpSfXoyvVtlA92qAMNzDrCPiI5aFjo/sK+CpwMwU5qnDeUQu
QgKy+iDG51L5OZh1hYzGxkX7dBA/G/vYalUB1mphIntqfr2bubTZXosfLNJG25dE
lEcqsrCm2G9VMyjWwrj9PigQvoqt6jUtkGn+1FKEkxGEUapgKvBKfPYvnWA6f63M
zDuPP9Wkm8J9TKJj/NC6GHsu/FVbjqTAGW55ALNPBlL5FGnNEp0F1VkBVBywZ8eP
pszYLcuj5tnEcF5CGYN9q0NP4Ai9K7QAI3hH6b21SInkWgmmutQQv5fP9uH9XJ6B
3wWG1AefilPbCg3y+JVYURaKSTb0bpRuMS+FP81KW8SPB8g3mvnRiJAMzWZkNpd3
KtOmnF1Fu/AxbYbSnjR6OqlGft80vrHHgitfk6Ebx6IivSN/IY+e4LOegR7ic01U
EKJ6S4cxy61cbkeoGLVXY5SuqyuJ1KRD2qdjUTdjnUL8aXfFxwhXlLr7XuTAYsKz
6EkTLQ6T/NkebYbFwQHSi6+Q+n6jK5o1ohGL7ZM/SIWdJCfqtD5yQ5iuIUYu8+fo
WXmRlesAZrCimnwHFhrgicFgP6nwEkuvK/sIh21PHq29iIJ3+mBP3G4KXk1hJ8oQ
z+fYkun3OoiUKh56XVQMmcnYZI3OO0JQLsOu/zqEbrklRNKcIaUtMOcZhouKvqmS
V0oqvbO4R8pR2WLge+Mx2qU3Jbd6+z7DbzNwTSCt+qbXHXKnIDy/BqbhsnuOK96q
QcEQLsfhtWecOwypBIh5AirYSsIEbhHimHW4R0GV+KUt0f4T6K/zUDquPlkIEhJ0
jIs+kyw4TFMASrAngeZMOCJ0pmU3muSjMQ23yoD5wW8HIqqryhkyWOMzDnhmJ16J
BDEdGux+y7/Ed9JdZWzhQnegl9bORWM3t9McwC+9s8+j1iWnO0UFLfgzwBIH1D36
cBKOmDs2FTjtmQU4+mFSDg8+qKr9AkuYyTqxU+MeaezlVu7tjbRBjt3HQHsoqbkg
SJlU6354yScMSpQ/Gy1+Krs3VYLWIwVF36+5iT/MgE2WCvYBjXR+/ugEGXvUdajk
PMMYCDtoGQB6AOf8UsdR0Eck27g8G2wwocBNqD7Qpgho+e3s7ACyHa5nTxDrxLVM
a2rCi11xHNmXHszKewx+QRMKz0dwiUBnZ4doMxpxTxpHTuU/yKXbmSbKmm1T35Xu
u4ZAbs6L2EXJMzSOIsXEkO8EcV655ZGWZayM1DHxp3pgeJMye546g3Yxw0XOZ+z1
+MnPLtILsc0e56o26m85uRewHsFaH+dJNrQH2VkELPwY3Ef2BsQU5eKzTLz8cjDc
OqhyejMytJx03AHqBxY8U1MZe9EDBeg4sJ+elf9S2RR1fuYw55gN3LoNOeDEyqWd
l2rysrsKx2v5F2u2xL9exEIei3HssxmiLxD1X2XrMsAYOIqTJVxCpVYuai6n2CHv
M+HMoYc2KQBjTzlnltSwmMBqz7SSnok5NL18t8oH8gUwKl0X1UyVvys5GIAZDqeT
SC0OPt3mV5ynoshEEj/MPRDbMIgHl7RwZnlU+rS0gccOZDSPXrKJyFR2+5nDbhcY
EtbJeo2iNe5pCQjmOsWPqdE+mv9UPRZFfeWtpQYeeKQ9YScBUiWy/2xf3BC5BF4x
Q2JchdywiiyKftL7Ut4EiXJq0HPd0U06zU31oNygAdsO698wkrLM1BjvYliWdrM7
X6q6LI9dbWVXExyGb3iIoLt6CwAD+LZggdoBxGWHJJ7vlgYv3yE3+69kHZz7M3k6
yRADzixar4V8oNoInr42up29+6rOh3MYR0sS8nNRxfNhpnKm497yFFmX3MbE4IwH
RUMp5QYCz3c7NIamv4toXQcnNl8nZUZspBVPAoQdfGUv6d1QV+t6ti7jkU0Szv8e
uJOLQ9GIRgYoSrpYBNWalGUQTrLSzq5de07X5VawBskuu8uqBhP/nak/NbJHUdZH
JAsWFctQW1Telmx98JpXpRLXodOxfVH8T0rJNjyDC5bVipTnU7wPZaBVO0DJ/ZY/
l6Jid8HXlXkwfk0C/5Ws4PVqx0tub4cZPKXCVJLPcvs68HnHZbgTGsXk8dXNIijo
wK2GvwYa+XH6FXyMKBHj1G/6Iykghgs568TK5PeDmtAUhvWqWsFUkHGEomeTJYG3
bWS63iaxF7wGSMl4GSahlhBYvCmpZ0lJwOm4PzeeTURxrrdBZVE78alSWTZnHwMH
pNL0TMCunstWnSjZkkknSPJqqiiVSSg9Ox9mn4KJXtzzfTpNWGKk5XACThy8DbSr
xfL1EiOPcchQGWTN+tRlZm5UiN0BtWQOpEYhj8Rh3dYaf58T58zAyjISZyqdJwI4
um6nhCqKvJU6Y6S7K+IEzgkZ+uBtntIAf+99SgPrpDlLP5HI2Wk0zryLprYr2zRp
GZGcsdmRVSvv7A/DrRTjIVYYWg+0q/5Lu2IlCdzTI2YZHilpmyZkLsvHYQtjw3QL
bJLpuT1A/A0VxghIrWQVmNzb71sKZNdfOEuw73jNCq3cWDTxt9faprKx2DtvX4Jw
WxM2bUAbLmgL9FjHhw8AJRxMA39caz30mdpZZqkFQahL/TEbUV2y7wTEnQCifK0A
yJLMC5kqYCpoEEjQX9T8+n9sLNqIe55Cl4/OnQydsXcujZcrFLO8C5Me8JZK3Qmj
YihvNLwN3CheSuE/JQ1I926ckikjdYFNMfWIWTDwZnVqE5oRfuc1CB58tSH+NZrR
olZhBXubskb9lLpvz/DsRxXCXzl15QJPaxO6dHHo/ZXYN+wzDQlb9n7yQnyVG/Al
oySsWbl0Y3dzY47dNeWsmFRG5ApeNMBwOZP5tvlQbue+sU2RimOXngyyM4TrBvPu
zlqYBt9nU+lQUHhbfcUj7/c3BoCCb4ueixy4vuRD3XJp3zXN4Y1GnZnM9a79yq+o
De0+GO9/mWY6aZOy15g6ZqjP0UiNih1Vx0I3xFGaqqOjw3xTP9ESD0j3dLzthOJH
Y9eKdXPN5NlV8i5eRQw4YilcgltE0B1h9gpKb0kfljg2+OdaCKYTonvE4iWaeh+1
m69qTZxYaTSxeYC5KxfOEyv9x4J6e2FFfRJvpyQcFMHunMDCFg+I0bHTSgvYK5Gs
6+fKYrQzd4O3x1GOI4BG5IGwk4/zUrfQsYtqkQSsNDIuPVVSk+8CXIRnt9TfASxG
GjgDBjLkA78mgRoHVtKh2ziyA4RLzisDSLR4EQfAcUn4Qj6BaDn2h++RRmrGWogw
bmCjOvu/5LeubjxxFKA/HXNUHrwI94F4r4rhwmvQxVqrCSs8JvZIol79Q/HfLA7Y
0yHU5nh1zEAMkriBP1zYNAEjNoiH20NkkGwZszWjqEZdlQSGV3G1s4dpSfw6CNUs
K5FpGbw1RUh6SAeeUiA+b7Rk8zdqmxx/80Zr4rFP5Ys09Vn0JBGK17a8sI3Gxpw0
MUHHXVp6dN21hY9Mv6UKYcpAcCaptX7njO0zYxI4nHwacsIZ1i/Xy7VYCyzfK+nO
VNorgCx8weJ3w6RlJEKM/K+RrrHZJcWaMV3UfQ7dmilsdLZnWgqLNBiw0cTUPZ+R
2B31z/KE6MJOkUV+XO7/qN6qN1VWWOUAOduoCf/bvP6wLWY9fbPZqRprxutLAt1x
47vf1z1Z/oTXEZqiw5DWTVsKPnRPKZRyowK4Ei6PObmwxq9qSnVCzwcKMIKYp7QV
7i8GIMDr+gpuKxfN8fhANKkF0uXzZScWpoRfewLUw8F4IHss/hnCz61DKcv7Km4i
d2f7VlIHjoaApmWiUjmmxVDz/V78+NaD+HZtILiJAz6fFK8HZcQ8McZDFl2E7Ugz
VLXiCemKXqCEzztUHqhxckFd53fr3bVV/sqNIF4TReKLGjNnCj9uMC1Aw2WjC24O
FuQR0n1k5uTVbB9EBO1T270dPX7th69AnI/UMg+YVOk4G7HWrhb6X4FRW0OlsNOk
sAw480onxVNjZbY0CiJVPzIo6AdUGQeHYO9ruefZcJMSn/TwBLoFaDumfwxLqRjg
vZi0OUqNGe7RM5Qg6xJSgaqmaFc1mkK/7nzK+dNk+qpWQSwy65H14RehLiF7CIw7
9ZwvmcJNrnxqMCosdG8hzROCAczBKrEQBlaohAew+PI4kHX2f7hcU+aTY/p0mmyJ
neH8xTlOFr6oR4Lrg8pN+Wgsr6MC9QHEb+j82AaHzDPsVBOQq+X9NzQDe76jtO6u
Vt0fB6S4QmpjJ6CLGUG5flHuMRf+KDLAt4j+U3TuQFEMd5cCidg4i1ACtbs+qEef
J+tUAj2wKZcVjbNGObfi0XYu9tI0dU2+12HNjdUf5jA5Nzlht/baLv0fPJaTGcS6
wvxPB2ZoVcTbm+kud5pAEkEWWRZ/e3S6Kl/BVo4kYT4NVxnBvYfWGJ8RNC1lodbK
KoUqthwbrx4dUdV6K3pkO9BW5HWLZkx18oftoLvh1epOjoHPs+0IBnl7kLa5pbP9
XmD4Q4DcVc2bEL1aofaBJSgjXHkfAxiB7Wdim1mUYUac1Lh/nyYtHSbLjXFkkcQh
ZFk36BiOBzo1Jx6n0omUEqkCEuXIZ08G7GLXaYiDnRjQYlA7Rx1kwT+rtdmy6zhe
Eiwho6wpRW2mxOMtyIy+Ux9rWTkj5z8kSwNmsacYYobKHM6HnenM5ITFYX7Bpt+V
0IiozIXIV7Ulvg/hlTfqSXqPllE8Ct0Y+EoA6AJXUlLWIGm/eHFKFAfeeBJAY2R7
VTV/hUu7O0crSweXGGSu7Tmw3g1L49idvh4uNk+UJb7c2Gyb/tE86dU2Nrlc7DWK
ruXd0GxWtTGU10f18J/iP+55regNlGIWiYMPbjo7vHH3gDldh6+AHPfiFr5TQOmo
m6T3qdgbJ/mRe4xqoBc9XhVM8CxePWG0CINEHCFgGZbOzvGy69py7dKFuRX6EfwU
octFME4EPaQ4nQMRxITIyjQ9RiMQSwJk+LNVM7PqSmJZWolfdY1ekTq4ZCUiotE5
dcG0E8HfWRUFKPIybPITrEArYzj5zB2zrXvKv8MCIJVXdmb51C/JtB7r2gQwtqyl
m2oFDVcdbsw7zeIbiq9obZ5srIhWa++LksXZgbigOZoqvgxrNUFoAvlTLyOwRjN5
U4Jsr/DyYuIw2eJgc0wnmtf6NQho12TD0bdFAo6c/hylCA0EgYWBhYyV3VZRcg6p
hP641IzxnsGZB2CLbpvtuVpe+r+J/ymZjDfbvWkn2Bw7K0ggoXCrbjKPQ4qQQnUS
yHFFK3YUk66RHn1gUCE+ftsGfft45suR3T8ZtPnCFYIHKhNwcHVPXf+EzSXpRmho
HNs5q8Spm32QkqNGXMy8BsQYPZKHhJmtYjZ75eYZbrfmA6Z5ZgNWvZnLuOU24DIG
CQGSGZL8TG1GeMGyiYR3ghusEFni682So3BOdE0c4tGHluhIDi/2ruqiuG7w3Y+h
wIwFCUXbNAPcqpVkD4cCay61pflMgq8NmIhUH7gptbKKMdvOJCyHmJjb2TZNr4RF
yXcNWj0aLK5sXGa63yJ8N/elPLMgYxuNA7x0RWykjzrtU5amhMy4q04jdvuHmiYY
IO8nRDroF+Sp9xAxsIYObXNZ/8eWJi4T//vqwz0DNbES7CIN2gCxBQYRnJrpM7XZ
+sReDCayKI3jEoQyVDRCBpgo9I3Y+YCRwwdtxGWm7pqtv/OD/1ko3LF/KWluRgna
kkQ+wTjDBeL4DVFVtIoV9c+jRgbFND3gYLpzFJTzHzPRS1NRQnu002clDn2r4NrO
C367gJlea1WTZ723AGU9ImVwHyJmy65fPVgGMdT8TbzMmRqvcZWxPcbeRJgu5/u1
RGvBUBpB2/NFdWGY7Zk+3BqHkvJ77gl2/4UBxUb188zzukvRqCvZis6acdMSfWNK
i/lVH0WzDJ+pkfje3qOBktK85LWtgp0V5A8wbpCGV/TaUn6R2JQI1dItmNNvGf82
pgq0AAf4ooT1rgaEN+AoF7W2K2/ewh5o1bwTbLYbw6W4qq1xEMrPf1BF5gQHB63v
siK5DWAqHTO9S4qu/KG73YNwwRzs2xYQNRfab1DoM7qZuPO3FACl4yFJkQrOzPkI
g9K+gOkcy4ZvrAg60pGZbztW+eZGPVOBLNDMmjmywAKLCX3R6l6VH/BQ3LWE/YTb
HuOiOk3vWOrfMRF5IzT5tnVvOj+REcwawAhr3rpMmRXlLxubBaX90W5QrKfLcSNF
Eg6ywWRW9FNnDCSmYx3BDU8Vn6nLr+OKdiiVMU4pk/Y48WcA0opKEjl63V5czp25
CQufrSd4bleMUxSIMJK0fAdGcuMVjDMGpUkES8ZaTfKTRRK+mEo4Vaa4k/gU9X3g
zWjOHSfez1WX6TlWDWLOmJ+UkpzlsVIBeIRFF0rMxNFI6l4id4phfu16zRDmXRM2
zLNGpGmilKLKZuRPiM5MHru2uSPaAMeHYfTcqIAyeZkrGF3bLEmxAWfh/Pe4q8Bd
+GdPBNvsoIDOKg/ivEsPlnZSSIsu+8ugW54nqFrv1Mhct476Vv1onPRQXvsRYn0E
0ycKGHqRQauC0Q9XAR85YgHf8els75Qyg1S5w5MtWymRPogjXahubd+bLx+HuXcl
8/90yTc8L/cVGmMJgInUk4rwECaHh5geeL3SQzpYGPCd17DKWnVVW4i3jBNb0VL/
+4UZvPA2pIpMx/az8JJ8KQlzF330yufUMR8WpBmnyzUZqsUERHvAGgHpR5oPT5NU
8AWkiJzg7LP/8ZSc4RI0/YQjQw2FEXanW3hGU20Ac0DbHD8mu87pcpz6+qRxRbDQ
f07RoqL4qcv75IXVprm4Ndad0JksXyO8xzq2oqzITzsQYYYhlYJV6kPqM4NfrlKC
mF0d41ArW0cNssFbUV6pyPGGgJsjuTf/bJ4XoOIh9PfpwotXe28AT4SqBFIIFXrX
uFxP5X6dYFlHIq3iADv2g7BxlNmgJWKfO2YbU+R1CpgVFrKUzmF2UxenZFL8tPx0
Zoq32+ndvU7sYXFDyECS9ylOeC4FXLxjnP4ivABw4kbCOnqbtcBHJ4fZuS5KzD/F
5/Wqxqel0+y4/Og35ZjL3UtjPj5Td3w46781bhro+THG7PfuDdbmQvhgwN1FvQAu
pB0+UCrFKhBb7chvzaa3i7ZucfA0vThKH0KNoYqGAUfDHv7mMXsa98dFFiD5NIen
NibYmPGEXFjscxCBPS+0TPsBI4MLTL3zEnB7XCajfAWtipRZdCkZmjwTmiOFp8Rw
gHGwCp99aVFzIqv0o4yN/g0uVLcy3vSBc5jDjGY8pmZohpnFLNBilTzrRaCk2ydn
t0R/gR+C7HJ9Dhb/ajAuqGp3ZfkzDEHGVZXfWk52/xluazySNbNmvcEr/oyNUYhL
mDiG8fzjNyFNuzor7YrMC7aa5mescgum1hsIvHRIf4w2Q390uA3jJPOYaoNBba4d
MHsBjNIu8hZ220PVb1MhMaPyG3kUaLgPc71ASHSK1j/elbKVnWDxxmzeJ5URU0fd
YMGp2ZFowUKLcaQ8qKz+GpmtnQILevoFiVE5JiiH0Zd1AQSD9HedogkCGfg+KkLh
U/5Fxd/L3koZ+IqotTu1+sn3lT+psMNzkugrp5P+SFJBkYBXCpXiLnbnKMNxYyED
7tk7dYI3HY+ud9MfV7fBvcCvde1tvo38z5M4NxJ0wU7mfQKYdKOFG3kkYc+bJizj
fgd+2Z4V2hqeIdFKViWMQg+ZvagxlsS24/FHLMuLBoT1zxnZqAGByjJjZmWEPX/+
/PGAnmIjtkmQ3/p/aT+EklL4lqMJae7WxiQHz4CLLAXfiKAzrGCaC3pnYpYD4MJw
ZMZo8H/8EVPj4ZjPu8bDumb43b7Dzq0l2uLzexcK+hcFZrUxA3sGvpOiPYosragF
ccV1Kvyghj3eKKFa1y4oB+FGkokn4hukRpHZBvs+glsaTDcpfCrrMi+e3LBRbLHP
QYrpYK0OeOD93hbIWJ5iMHeMnqwKahX1AIA5ixiARqZRHQnI8GyRwCvWt4s/ov29
Nb251xYqRIW+MBnEuoMGiRPjsVfMYl8WIdUUTvGpvsujQdg+ZTyMWNgUGKSAE5+C
tOnu8vih2TIOg6II09zxSdp2FAPYColQ0prciB83O/6uVCfTyayioZfEZS8yBu7k
oCvsXh2d9NsNjwScQgjg95ZrGYp2VgZ8N2E3P4+14bBVabG2NdoHy97KTCuZMu+7
5antChIKfOYrLvzA6A3067z371PkvM/M94Hl78d7BRGK6NZyEqHNH0cSl3+SIBqG
wpc2lxIBmN3eVYV84UOYW53sy4JIEikWVoY/BNJjAv9YvhyqOeZ4EiUtJ2RL1YUo
MyP2+FEi/+dAHhmV6nyyJUD4AvueEb1YedkhUXuCWbMAP9H3L1aDPOLOIH/458dr
KtW09d2LLlOf6JAXa/vy0TYg+rBaXNzxSSFqKVwddpB9s1PJjWuVWLr3qBvjVswe
xl4YxSjR2ReF1AmA0UlyJtYqlZqwLKt6NU+5WEp3Mq/ZQwYThTSDG6m2YL2IwYQz
x0rbl9FWdmdFyAYpBddBsje+2gPxHkgYBXJW0ks78UI8fNFjC/jQChqf8g91spZY
Uu7BtOjf3GYcGNkBdCgkeliqBQpD23WDF/CgLShFM8AKVVQwQNzdFdaD6CrdneUY
7r+TmcH0UvloR/xskqoIs9WwB3tGPwL87JaQreaa4wGQJR3HEG7scGO4z/nbBg07
vuyf03/gg2lK3JISnbwE1h9ULaRoxOlJEezFkR6CE6Aq6zkfXErzFQF+NpxFS5M+
s0KGhibpsDuB2KUDNG+lwYCHckt21fh851chbzoN5xY/S3oTuS8FtwHgBxDvBUyI
UcOzJ2fBn01JGha+YB2PHGO5A6ZBGXHs7Lzzmxo4WJDgNmOVfJpVBpmKPc5pqMZ4
Rl+q1dcMMr1Hp31brQ6NYqwJtte9QvYbHB1JWVsb4vX1UUO3HYB55hptmz+SZ9oU
sSd9lVo+N96TxKo1FZ6yJGDC3IZ5a3QVmiMQA5U2PHwxDVSghEuVDtdWDjwLh1BC
vWMdZD+q/6z46+pEHvZpFa08EY7DS/xmw2zDQdeOeCol1gcKNEROlkdh/D+IU30x
L8ASyCOnQHpnHO+h0BIQi4j4pqnlZYVPmWN9AxcBJjZRKvR5rDLCWg9olcqTP7lx
urxSdJRIVfI9Vt/LeFNOJustMT4Khc++8VXZ3ay8Zz6E3k4o5hEb6JoZXqA91+OG
xPHzxSRq6jiHI1i3gpJa4o1IeQlDkI71/VubDxRTMYdyx+n55jqBWIFA3Nwtymln
iD1H5Qpt74BfLlFGI0GYEZj+ruDFdNQjkCPwbPjhcySaEhpajhU85LQjfK31Bvou
GGSNhoOwfOneWqKKzTti/NZ28PVdkom4qgiJoUNnYnQ=
`pragma protect end_protected

`endif // `ifndef _VF_XVIP_DATA_SV_


