//----------------------------------------------------------------------
/**
 * @file vf_scn_gen.sv
 * @brief Defines VF scenario generator base class.
 */
/*
 * Copyright (C) 2010-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_SCN_GEN_SV_
`define _VF_SCN_GEN_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
E4FsF7tweV3u+3S5qW5bvJfd4m3RguxlL+VeaTVUR7J83INPjSpNqr+ARlOnsfdO
Qd0ln7ZtIxyKaWLVYnldX16g2vRQdqqcjDN647cBMzmVzfaFR2WA6v926gHZi1a0
mwbGJScvIswS/dxCxK6E2qnZ+YTxUpVGRuqkUniAGqN5YSAbLP+0+0+gF5F1F+Z7
mJGU95EIOcgE1gijXWHB8G3vix/+uUQCKPBsp7gh0+NC56YqUuEIQrHQhxf0QiqT
s7bGsvLS8MOCn7Xi654UC0eHU7c0+5G1YwzIw1dNotR+BrpWx+dEmFOuerESxtT+
sTa4aP8JQ+XFuGuCpCvnoQ==
`pragma protect data_block
6wca90gEk1BzDCCKOOMtWd6WOvyS4IvGlCqC25DFzjNoKd0F9zh1hBuEit68wN/n
wp5JmDrW97rMsk/2LjVi6tBk0ja2eZsbuzeP/dHyRzLyy7YKqnR4hmwb3RL1hWyB
23+uDqvHrgnnw6WdJQscZIAyKgjEIB6Bog5aamMFBSGn3ogbPMqKBX+d48WRwCUa
asWwk/S5VoUEqFNJCRWQT6jTn/As8lL+tB1vKZN98gI8w60KQBFlY0HE0rkVeVk+
SVnL79N6VfxyuhiNA4F6UgO14EJc89ElU8KDH8lK/Mhv9WR6Y1je06ypcf+4t0+J
vzK9UFOYDPVvSfWX/Il9weqP0fGxkf8UVKRx86smY5yCC4V0lhu9ljG7OBvKAmRC
5q49Yo6nmJjur1qvuRNklyoFhcKX6cEzGUo2gge/uum7IyAYCHW2RjgxxARU8T72
1RLcr9dEroP6A4CIfq6x5fcfMyqZSiyGPlAjrkN0cQKnXcLzpUDXAmiMKX27i1UQ
xzQO3Ck1ObxWUQ9/jP4a//6iJ6YWe50SQN3K3zJHepsYAt0+HvFC5WEP67EiNw2S
wRh9V4msn4FJyfVbxjXzbL+8joBZdHFF15GyEmUkm91u3jlUG55yhTzTWAppPOyU
eRo2Z45LEpNwzGgY1hoUrLvg4BsOIc+xfxfz2WG3RuIjdDZ8Jk/rbYcjJQtSUg4V
VOKI89j3Jib+hQ0KwttIEeJZc6udSb8ZypcfthWFRArmWPPn2ca3s/ILdWtGGHUC
HFHjfjbvvy4XA95vs8ji/7l+Zu94G7Jju34KiYCCWBYlfeIaeuVgQO798B28YJDT
aVUYw3hVNArFgHAh9/vJFc466fLEY6asjfLbIZEze61PhVbqlFIZZdIGS68N8Myp
p57QwpI7uchgNRwRexAWMOWuZ8e45dpT3eVM882axlv1L/cXvA7XaDjpUCY/2CnG
xpimV+nvZD/GRfxDKBz4yu9je/UPdAjqSFzA1fm7eKDVqWvRs68tV2AhRxHCaaDd
2kQUlA36xAkMCEnM4NZlpvhC701C3NwViOddPgOorgmPmacRYN1ktF54EFumS8hW
06P5dQqEXXAVy1qR6t6Hv/ZhiQXY8wBAlV4QNXXOdlcM0D791on0IeOtAmHupOI2
532LcMXxqQaehdJipKb8SOODW31tVpWAZJjyNk9x9OFxQurgfxRwYxLCxd2kXnLK
I0f2alzV5iUCGUviqqRrkNbVjoWxDs2hzd5nGWJoprAE3gLYayeaX3ZkO99b48T3
EybbnIFV0Vpnrrcw1zT3/GP8NPxmJAqQ+OBO3dWXIak385KXb2dzu4SW4lsEPwlo
xUWEUoOWCrJgUljziC4p0ItMgw2V+bm+2zU0VbH1zRsv9wum6fD08nJycjmGOZ0h
mYZjO4l13BKZlE8/c7dj524m4rvZ0Uv48D+hjn+cerz9XN8/HockeDihfk8q9MXx
XqWyBVGHmC2JEIjBfcWyXuZs0a0rbZqDsDLFxNEYUs+I6DV7isM9K1W8NiR5kDFT
Po7SO7HvNsfo8I5iZgAbYcHqUCNDDSkjorEOT34Itz+IA6gwjxbDjhCNs7WuSWdA
0EyM715r9apJqg0/eBaSGGxudwa+9yXj/sw3CGxHISsHLjmZyQbyPnGNP9qeAdHO
IkOxuQExhJW079WrekxX3U+2Kv69E+RpStJjFn1qSslouYoZmqbCl7PrSUVPXzLJ
K/FcQ9yU5cgUm5S2LCh5jmdO3g8C4tL5uqsqxviYS82zI+lWNmu3OYRFNcC4ndFC
zws1PqlRVLxYlyQzv5PIk2VPDHJGgzXpu/iyZ8nIqE3vSwjzzN3Y77iTXg+wWdFa
FWuhMpupN8Xa3gFyYazv29ewvVIfT8Gv/teOe7/R4u3cKW+dsZ/C5fS/atFEe1sv
ilM32Sxdw0x4fZfz6Otd0OEvETdEMKFgTbINc9Gopropzs3CA4NCNC1VQc0rl7Tk
GDDkkrFzGM/6uywcx7vvNVN2Da7o4K6hdTgo5V+ak3OtvGGJderIttfgWlZhCsJi
INmpEPzSY2dNLVzZ2kvQ+tpQznrCekNfvEPVEDVLJtDqhiRtZHjYlgkrTBWpJFqm
OV1Y+VScFjGU9qt81lGNcle/W0oB1zGuiOyuya1YrLGxRV/9HQEApAtM0G/NCgcL
vq4RIgKN6ZEgbsow2fviJKAHCUrTSgI6NRZlWoFtLjpTz6EvwBTGcGDGOrD08Icb
9fNzs5JqZlxNHq6n04L5WaZreaSjELycLbe2JehPh6yVrJTNVApwXvliAlfTPY+3
4FXlyfcTV4tvVFvpWD8t3ZukQImLloAx1zElxrzWepajUILsWTQu3lQjfWPpaGYx
ezB5cdc6JqhfmiPWdRnGRcwsl/3LxfZ7emLEkvkLiYOqYsQJx6k9X8pnAQdUeDOX
M8kmANbEg3MueLiulKbssbvAKhZTO3r8qsGG0St84vR669a2+jx3N8qHBl+psqT2
IoOrA7O3oaV/Ql9XKK0ft9wSrif6lWNK2MHkwG3y0Qlnt0A/Zet05Gmr/FFA8tOb
GO/VCGgcNhdjtbp6Ae3SPuiB1I4OGk8/LNXcRO2RyXP/WM5yapEAMA/7Bgn9Idkq
r+pl/FW21i3eImw/wGg3rZXj8Laco7dLZKa5xqxMk36ZLSR8KipDdtKOJHPqIwJ3
xxjYSIu0Q4mEJ9dArSOB6eb5sGs3HRnD7r3ocvF8zEtsZGSxc2eafeQS2pSPs6nt
LJfZfE9t7GqCvF5QFePHIInCu4g8hb0jvUu5x3Vdz/4V5Cpzu3vthBm2ZkVQv9av
AsvZ2SM1D748O2/fkKhINdpiXL6o+nvZSyM7Cd/U3mR7y2tk/sqyx4Ei3E8tXPqu
l0D5yzbYpB2I/xL5PnZuVDh0iMF3eEYXyfqmhsnPbjy91T1Y1FzqzsjNXX23MKcu
quVZ3TDKB6AD2wGWNxg0YPi5i8pkKg/MSrLJUJav5J91Tgi5JFpkdOMPchq0Y5Pb
PfhPZfMoXXSZxlQwqX/QLf7vbivC+OcoQ+8xsATpQg2B+vbiZIo3u3pK6xSLDhC7
QPtc6j2greYCAHb0J9ZmcVd2LJ0xAZvfYgHIlAnijHVSzKGe0vvKgmgO2+/jaLYl
aN73tb29rL4wCtqQI7eORxkI5yHObfInyN7QnSmPTYuqwGWN6Q1u7p2QECyx23Bl
Phq7Llv1j3VzaXiGEO09LwOQnPo+Gfi5G8vDrYwShym3quw+BT5vSWXgrWfAtKqs
ydiIrlyvmPBcN1EEi2JGAVJMm/Y6NZM1M6HUG+NXo5jJq/G+bQfhF292AtSXBXsW
OIcPt0WVZRBWDqd9a7B9DIOz2WFvlffKav+wW9LFyFQRibeTz4hLQ96OXwaxOdkY
6sPtO0Eh/JRfPs9YaRXmWbZwjskhRU00tb+oRzJdHc6nox8Swg6NBwEEKQ/xSoa3
zn5q8YXhtEsZLd6RneB+i8k2bkgNJ0F2OEuueoZdZEtzY+dC9SF9ChCjOXGLsJ/+
qDvrpUsM0DhSKUEQX+83Ey7KI5dMZZLJSS9i0k/xmA0OrBWBciQaKdahe2DGTYzF
dWfked0LVDr2RoVlKEUiXagLO54seLC0yl7w53d5hK9Rd9bcumZmP4+J/3c37VQj
nktJceOhoDuSWQG4rDLE6nm99o7CDSDx6NniMjaDDQ+eym/TGn+fPMMp/e5ofn76
BuRgp/G6YvfPf6tB3oTaHzmiFe8BnQYpBgovxvWnKlV9djF+JKR7F9suC4vEZJkI
LNhFTAUGuw7mh60mXpbG5OA1TdOrsNMQw05hxhcbKbzHEJyoS/1CzQ73zLwVJL/q
0sRGZl3Lx88LO7dWWBeOBtbMbIRmLUWeKVZDIbJR5aaovYfxIcSWQ4sKFBGH7vvI
AmC0O+GbtrSTFZ5gZygLqWIO84SNMkAOV9/3WaNv+n5UGqFtdYFyivBj23DpXsKP
r4tRuCjE6/OkJ2oi0xEHXvR6rEraHs6ya1Qx5cSRfcnDW/6+tr39weO/PhEsCYwk
BDdYqqbRLdH50kXpNHCkjQtFLvgxwWEkYqmGDRgrDtxl+2pMyzP4oSq8TkBApg9X
r/A/DY8fDVLutkSnYgIKFZFJoiEuw06cFG9Y61/UWnzJAPuMJ47w0KK9Oo55oTLZ
hdmLyuPkfewtgbvBeYJQ/Hcqw9L85cR0a1Vg/iuZqzIbM+xJ/YR1LC1mHzcG/jaw
9q2rpwLf7hR47SYUCo3zwPguZirupaGpsESVEGHyxEIVdLqzcD/6kbSgm7i9jybJ
Vy5kni2ACR2rT2ZDO81k0WuaZEqyZHSYxRzirMN2FftKTYaKFtJ/rQ6Qs1PpwdrB
fMrfbBFjaCAxCn+9Tp82PmMPkEh0br0yuoDYsGxb/c78F+UbseVYTFN8+0I5E5cB
cPQzxuGl7z2p0yo0uWsGqIfNRtAEk6SKJON8HaVz8pszhp9PnMwgEb3mT2Fb9RMC
yhyNn9W5quRmQSWfjp7/Zl6xXZTIGFjzKT0ugBlWWfmtHXt4dmqnC3/Nfz6f4LGv
BO5cVeDeiZ8bnj7Bqx6WV+D5E8E9ZKbzfzjBu1oNIAVPZw3fBYpbShQ+5VEdgbqA
/dtMUBrfT2p5CXK/tAjH2lDH3qRZf5DKDjM9q/NxJh1OlSVUumgAxSTYHZ9EZm6+
RCywuO+m0wO8fMYVozQ1W8EqXWz1MJp/98tPMDP/DCxBr7/Jz3l883knuS+NU4Kq
El4wm4zUvKx3tnm50aLiwdVBjqoSyPJCPo6MMDKbcYBmRaKK/Y0W1/MNL8/chCj6
erRaUUhK87shTAjGZAslR+/HFmTjI9NH1JWcZE4sJsU3yWz3qsQxMobvK/ZPtIfp
0OsjNuAjs4EFiFboD6YFES5ocCEZiPuQbOdA87GPZKh9KCDI5YjIL6xK3u2FBOGv
+0bJX6m+py25vyiG7wwg3lKBuTefQpODvpz6XKUcMKx3GHRC9tDx/8Fg//sqWkfM
G3dfVTVQ5Qq4w6EjH0cYVD4L0tdLO0fHOwRHtdp/bBxK9driOw0h6N6TDmpWXgXo
EykYXKBYqkPsra77b5aX7X4A9PI3M4PXAYnz0AdiTAEJIatFqTzaGVvWDeNqLiWl
JZpP4TXhtcxTkPhk5y3BXZbg+tBBff8/9DrMBq7+BdOaF3y2rZaBaLNnoTnBKJGP
6kFDlAd5Hqo6D0kb8wGt9Nz6Ofz/WuKEGQ5MmU6aoNWFDhz2jF7XlSMZzWV5VeyW
j9UexJOUNsL54ycq6bzFH3cgc2oI6u7rzNowvgpYIFVcmK3y8Ddp3zKyw8U8oqBC
BRcdBf1WBWPa/lSpIJIiUjvHsLMQU6I6+JODd0n+F530qtkWqi0WpjolDErp4vC6
URtgI2KChNrBHa5px+zSHtHkGERmTKr5Z1C+dW2YWutbwjuG6I1ccLQw+UPGVZby
LirW4GS8+mMPcdFv4mWomO4EGvXnnPftNp3qloOcjY4ZmTlU6wEFVnn+CtaDQRBN
ajLV3YUTSUuKY2JSmZ+S1ygBIbQOFyo10oQx/Ag5GHDaeAhPDG1h6OB3aVRSmPfJ
iAuLtXiQddEo7zCCrmaPUAnEaFC4B3Gmvi0lEpjRwVgdsLvdH+4s507gbwGD9NJ7
hC8Ea6To7W2f1clNJTpxfpIdgd0Z31fbs+mZgmns0qpO3BRA+F2uXjNtb0pOTUEX
37U0Fgtigs253VJZzmHqF5ec/PlzAq8uZEZiDYOFyIfZJOzw70lJbqBt77bcqS2y
SzNg+hIHkfLClhd/PwvZ95sFUDRnOTuiJahfmNxdNI18dakma4rqSnkd2XKA/R+J
SxuiAg6LM2Qnwp7LCjUpaUqwxR+JnAZ2UXZqe+Dw5HK7qF8eQcN1D9iw8xxKZ8LT
0bKLkSLeoJcSnzuKg5W2reP3x3dDVbTYQGnjLzqekWBcUkRt72py/RQwH8xTu0p/
Ihd8714zvgrdOpDTrCQC5Jz1jQSNE8WmwirwZJy4xbat6QXoOT3NCfbZsqNOXvgA
gYQuHyNesad01lIn41axpJMfNGJrSzG/3j+KZPUzHGUt9HyNzP2r90EYqaJSo4R1
n9bZWn2AmJ4s6mfigx2vHAWknpNjUzZP7MGdBPBIiutzOtJMtjdrZ1fwVkiyKGhb
Qulf+C98jsqs1nmWKALHCH3lPYJY61TjB3mSofMkO1GKuo/1ldcqq4IfqFB3W7dP
IJk78SbwvL7lHew1qcgaPpTJz/OaXxzNKDHc54Mm3x2FTQZ81msNdEXGbCRgRtDi
4USqlcuuNNwXvPa20bJA7WKb9X+f3vKZvrhZBYJsJwMR2HRskRU6IjyEhrGTo+e8
GDByvqQoUJ5UujbO0n5yoF3XQ2By/5fYTBPt8Nlnf2r/G8hpF4uc3VbUbvyzUWY4
Lo6BKGjY9rEU9YbqGTtrvLSL8cDDtgpcbSPA1Lgtdssh8aohgyGwzCU2KyK/378p
y6llJ4gWLxMSPkTOXg+p97patkbb0MQ7waHXUmcTP29dtw8nI7sOsdZVG4DM3bEH
yTBnvS74fWyCBZb2JgkH7NLqOjAVWkC3MfV6786egLn79aRooLcO140a5KEIMDEE
Am5PlXBINer+RgzeBexHzcTe1NcFaaGGeCAft/RCYC2n6oUdiSLNULMS+/roXNOG
NmttQVsc4u6aSjNKeGCHBFVzA8FOS+2lwqLCgxJOc/ErfxqUxag90Yoep7oCUNDj
2as9pH+qqQUoCYHFKffOkon9nTyzDOLSR5JkbSFwAmRUgksGoBVvEIA8SUQmtaJ5
GAd0EBqHxGthTYQ8cmOuDhMkXJNH+I3SagbgrVqliueNbymFrpEKgp8weXjRNxcC
3rHubEJKkJaBnkLrE051W/Ly2md3SjFdTGdPyFslw7Lz9zkEAwl9rht4rsqToPEs
tEH1ygMFIAY5ISDhZsvvktv72M+dBTF38fvwI8qHXVMe0WkbAEA7aY0C42oiMm5K
jSPrYUPbEaazZ3BDf1nQX/6vBiC80HbZKZDjBeRB11zbpMpUVX0fMcn1Oc7MajDh
ouHmGy5fCjxuZmxQGv02HqzcPJtK2GA2k+Mmh0pYGrdsrriowmvVvH3IvzeWHT++
Hjg+UPM22DUHllTiUcbPh0RLwWdXkRd5s+zUqxgWXkq35taXesnBQIp/S2oR9Ubv
tG0dp9+/xGnKmcGzvRho78YAnpplWgg8eKJdXCnPbT+ugUywbVsWnkGhZbQNZgeO
W0whzZFYyC9YS7lb36nDMyBZyj7vD+84DoPnAarnU37S8OV+iq4fPzgEJNy26Cta
plMJlXdP9z047tv6GE7o412E4/hdE88G7A4Z8sWB50crkUYO8ORAYQl/4dA9ukAn
ZQKaDb9+XuAxbIcgioKxdwgXQlf3vpimhkSRq45YSP/5HxY2ODoQAQXO3kKW65Jf
WWQQX4XDRk/qHzEu1QakO90mK/ep/tGNWAyf3CAc80bYv7lpD+/iBYAZkRDEAOdb
9vbV7q1B10gpPTNaFAsh1GrcgOZH07crKS0eFSiAYhQCYRMRcJdD0gHYF2Xie/3C
qbQ6f12PCuqvylXAwMxvk4LxGbuFNQznGjz2S+VLBaHnyxRaeJMXU89QXmbR+l9C
iQ344JsS4GRQcLIYIUx/WjMtk57RB5t1zlszF8m8TZils2vqd/xnGXpqwWBDyr2u
IdXUxF7GnwL2TRBxy5kS5j7kWXKKnm17y9u9sfJMfzKihGYs9i0ouMu+S4GsgZXI
DzqCgwCByXSnTwY/mF222i4ettGfZGbrVDA6MfoJnxL10M5g1/fgCA5aLiyZFl0S
lRtv+QAE0rBG1/CQr67m8NMLhTdURDNgRb0/QrM5j1KGwSSiGjStskqtP6DIA441
lRYhWWchG9sgxheqLkK6M40ultitHbN9SPkm4fPdA88TNSiyDohASKfZdfqnV6p2
8ATRs+VZzqKTx/PPir2rd3nGaIDRxsldPLsAqicGQA7a0b4iXBASF5IEy86ODChh
UOkEwflkmg9rqd3uFz0jmWcjZMgn3cAzhPbunMswlQuwbQSrjkwuaAs7+ZNNK/54
ZgDQm1YRIAhorfbnr1B4WI+IMlXqRYxkmBoLBkU9z7pMwFQP24yluBi26aEtAzJR
ke+5+MbOcInCxghgtBoE//K7uEHjJ+b/zy47JdS0tsVcLRr/CdctCn6Et21GfLLS
U44/+mEy1XkLf/tlVRn/FxQ65Vt8sOwwib2DWXu0tNaXL7lJgNxx3c0Q+uAz9nCE
yxosYhA+I2GKsTMiZG3WzozBquqYK4IHJpgfS/nJAanAcDO4YCaxHEYGyQddhVog
j5w23pk/sTNq6SgqLwezajLEf0N9UEwd9HKGbb8BTAl5ZLZHrQrgtxa427r30Pgc
cBS72Bloca4QIYJTJBPwjoiorAoOZM4N4aziB61DrooufrFHd+fUNFXLzX6zeHzW
7ftnvpBTPSAFOY7npO+Gd5q0wrhwbIavTFA2/Xsc2fhlkub0X6AmubdcQ+IgLFXd
eHaVOSENAhdxfKeT4j45OA4mL80c1iJP9VajhJ6U13bm9veOZqTWPnDXEjSMp8Yy
+DJ/s/WJ2BDhG+/p1v+hGtbzv1q7C1cNr3lO2gFG5DJjtHYlFCmpzV/LNsn0rRsH
QSUqkSO2nBTKCpp2z+x56NjfCTSRqrowwKu9owD9asempBD1xKLISQWyy63HOVYr
f8sfY4tmtSthUezGwY49QpMJLZu5ClFu/fUCgqFHiR2JVDu+3nY10mic/YBpzluW
ED+C2XhIeAGBX2P6EQ4lu//DKvRjhESV2IQj4vsM4wzHXUtNRzR2j76iMsaTyPjs
GmQHvh4Vp9xCHauXkk8CIjhYXdS7zyBpP6u+honBbg8rJE6qQeOU1B8n95WLNljM
8v0wj38XYQqs4CeOyDQs5qDCWfndb1RTqMFxEeK8SV2HOPEdmTRfWDE2uFuSXu/7
Q8A/7HeKP4EddUTdJrR8OdoCuxCRgKdHGHT/A4VjF6S7wVD9bR+kHUrEcmZQcYyl
34xwnD98p1SDsU/DdbCPHUoeR2S8FZbjia2XeT5GhPUvbTzo69fxiIzCQ3F9QAzK
RFaq2XBmLp3lNOKq0AjX1tAei4+KQS/jubvnVwXMfaY2ADKZwcmy1Aye8Z3xBtOJ
LTmcks5qr7mL8EkA6LQL2ohljJQoDpjoPSKKdAEVnQ7RbMs5IjvaYdfXoAgN9lZj
lwlM+iP1YiNESsfaLMs/yx82al9k+LYvr1sTqtknvNypMZOUSKX8M7g0RqZm7+N1
yH45wBoIdTZEqE/IzGyqqjStWyWzZbbbCy4yblT55yLAGnRUQ/Ji+2tp67R30WOn
LjBIEo88kmgLKJDB7QetEUjVR9T8crwHckR/GKF7kte1Z5sTRqbJSS2M5Y8ywgvb
P0KyIbrEL0EecOIjRqUwHWeQr5ai6nbXcukIE7RrX0i63QilqetwRPKOBsekwqVb
668t4caQ3JBK6/5sVCFlCfiHBhh/bWccB0uIeZyYNMApy35n2KCDkAVC8IPP3+GM
Zd/dugE5CkfZdCWa2hMT4f0MLd7HqiG3/x8o+aR2c5h/2dFgb6uFRQjYt6azkxC0
oO/n5iT6yRuxEoIRHRZ7jt3v291sLkB9jrz/ItnwxyRzoQ5SPEpU8baUvRRd0ckK
n24TCEkV+Y255dsUQVHIdjFR1O5+LI5cg4J0aMNZIq1je0U0BWCgDyNcxr0ME1AJ
Kz4J07EXk99uvjbAfJH0reebXuoqEvihGkcS8SEPkq/Rc2kQIjjaRB2Y7Dgs9x19
Hc59H6NFm6qtl+wxbtE3MG6JTSq5ifVjCSR10PWAP+h9eyzpQmkKqL9ls8pjUEOg
pERZdhl66d3iv/7pL1sER2BHOAGU5IZpWIiphxHFtwkI6YNQMWn06G8SIZNPbd8Q
f3oOE75NLy0FtpEw3wIx8eVYX84l5YnsEt5a1AnbHsmsPZLi2SxSNk63YcmIekLq
qSY3coj3iz/4r7Z6a1RE1HV/uQ47gGwtAtNYB2kpWFmcFTsiIEMS5yZGZtFwkPyI
cFptqsiLyRJxBTPmm3wY8fyCZo+tZMlygrt3Giroh4+B80R6QlOkC4M+bvUBpUdK
IUDtN7NWlyLzeVg1q8y+RUlJ+CohZ3PYPGX5R6I4pS0fhv5aps5LOY2xeX96AIfL
i7rbeL4nH70cIPmEoI97eIlI8qY5GH5mAAcHlvvMqA81PENO0FildGRwo0BzUlh8
V1C9xp+xHLhmKZAGi82HgVi1IEOII86tSVEVRHhhDpq+XdEOh3ogDgOGszX0YPIy
1ONhIh6PopOkbBVOVzF3CGFDJCCh847O0POyfslyCR6m7SsbMRPnu3VTXCIJgYs4
NGpgZTtRtBdmPe9XiBnFkCJUU/+o0zMtkaQp4HaXDBbIocSvkuRNTlO3g1Aq3sxU
QiCLRTftLfArexbGc1oGjJWfnKV96WZIiUdYIfzz+Ig3qkTA4eLgGVHuWrzVzmCx
5bR5bfOzPfvvxYhcmoK7R5w6pAOL8aVSsAhAFAWU1vkMSpBRk81k5a8SmliQaZb/
l2ZbrZYikl8horPrHNRFMPNCcyMROWyQ5R9pow64HTI=
`pragma protect end_protected

`endif // `ifndef _VF_SCN_GEN_SV_


