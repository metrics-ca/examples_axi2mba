//----------------------------------------------------------------------
/**
 * @file vf_axi_typed.sv
 * @brief Defines VF AXI typed class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_TYPED_SV_
`define _VF_AXI_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
UwHLZrKQjRqDVSYWIMAIqlVTi8uja751X6xQRAg/mCX7/4BJ/qlK8z+Y4vNF/XL7
GGlzA2G8oaY1RF5mYP20BPvY9UVIpVLuMIC6lUadEN9V1knFeuUW5xSxM50KPZmp
qgfUKFVEltjE2rcyW7vDJfU5H5qTQDjXPVYivg0omrJELduigFtImp48A1Z3bVTk
RrTrLpi/Sk+b/Y/v70TlNG4RvbZ9dKd17J72ex7CEKi6rUQLFdAluHHjLOGRFVLS
QphsbrUH+h6aC2ZJ6AUIv9zBgYWQSZDOXuz7fle4ZTXBN0C3azbw0fPEBV+kV98X
IqRjGw3WUaS280UMRiTo/w==
`pragma protect data_block
Uvfnk+9vyffoOUWm1PP5gfAiu7GW4r0GvdU7fZQn5cK/TsArLGFoT0FgnT8tu5bs
ixZEvUy1MsEAXHbei52AGkg8J8eptP3AXlgXRCtKdxi6PdZYt32cf+fRfjf4dCC6
acK+zsnOi7bI9vIrh6Wm8hvLEck7QetdEwQ1yQh1haVN+zM5yWUMhmQkCingioCs
bMZ2HidWwvEB+su6YEkMPzw6txV1rD9Vr6lldlUFrhOYt2wfD5zLZVAOO5Au+5Kr
IY2HACKk5fPcV6DvS5VqajbAtjAk331ZbLqTdphq6xgC7fxuDHXwybNPPZn+ZPQn
UR3nqyQQzAAfwsheRcWzyEYEDjaOmOJQO0eXrhsouc+U1gKvkmr8giOWAMNKnLNy
8HZZdcP47y89wtJ+5OQzWGwssXcsIkD+bnz+koALo36BMUz0xVLSymWoR0AHoxET
OqddtYqo7Zs060mrm4Od7ToIsoHZQ5QTNj8LxxUILyeQs0gnuSgLjwU0SfVvYV1X
swYXdYFXpT6I0cy2MXXwAxWC4WAUU0ZLX9ruTgmsTq0xIVrsurPqKmkSw7PjakPs
j4sQce0C0jzqRLJg8ZWUOKA5WDlXaq6rhVfkmBe8GRRz4y8OhACVxiAyh4dhhan7
q3HCHt6OqA7gv5fXCTI5fDbo3ZbYtfzQNPMRA3kxcMBtvaThfmfNLULyctOqtTsc
8CJ0Y5xcJ7b5gsiPIb+45SrdvT8soPVGSJPL6ZuH/kBTb1Frj7IAW5hL3bhcWZ2B
GX0PwZYYwV4LcxYvaz/tvvRY1k76+/9Vzm12gy0SGo0zJYSeB0qVsQwGNK0gplew
EQx7ZUGgO0Iab/+4VKhAbXvxGCiF2Wtm5mdf9x95p1SIwn5Paqxq7/AeqhkOcBM8
SGDj1XRlzGMXI3FLymYoDdQOkpzbLwtihBmgabn6tf6Ijscij+L4nfiZO7is4o6b
+BHO5kJ/gOu1154OC4OzR2bPYjkLK51xwe+qZ/EfNWI8lXl1L8uXsQg4/+eNyKMl
sQGNraKZBuR4W8HBwdNNlyrdCUqC5612HaQ8MevQNJ5wzmxJgkuHOfZDIhKVenmV
FkFTrhOYdaZyAMuSFTYLxA==
`pragma protect end_protected

`endif // `ifndef _VF_AXI_TYPED_SV_


