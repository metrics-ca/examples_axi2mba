//----------------------------------------------------------------------
/**
 * @file vsl_sblite.sv
 * @brief Defines VSL Scoreboard-Lite class.
 *
 * This file contains the following VSL Scoreboard-Lite related classes.
 * - VSL Scoreboard-Lite class
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VSL_SBLITE_SV_
`define _VSL_SBLITE_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
aFvxaGdEVCJa18fRGdSgfVw1DBiDhJWBfNvkJVDgZj8qjeBKSH0EbwTBE1KuxHIR
sBjGMhAVzcKCO2lemWf/Y2QIYDI+8yD85Y+ZhDJ4gOLWAEFNDpDQTfh6vZde71YX
oraog3Tai+rORJPksawTj0E1DTxQFKbg6FZHA6JUrKicvN0/+wilXoCa+SALZM5R
JM9VuZqGPH3AE+OmrWC6B/fCSZQWKArSNk7g0ESCSQZ7Ctnv/89N+5v9miJOd5S4
f2+0yiFJsnl4Uox10eexVhnoWxEN7LaTi2e1LJNgO0K64IsD05Ht+l3uaeSpZsJF
G+3+8VkgH74dMyXCe2gQ+g==
`pragma protect data_block
kfN3cENJB4Y3aole+F/utNnu3YJShwxPp3Xfg8dRz75qU+GpcTEnixLq+VsSRPXi
oooRvgQDlYvdyiWwohWe3s3jIWfIB4LzvJ5GNcto4ZSljTt1nM319aMsek8xUSle
L0d7cnZjhPZ+WSMPsDRFGVp2nKENDuHyXSyLmi4E28XYiYP/wlvDlPLhiXLTU5vl
vKwACl2xmBb5LiZWZ6zzYkurAlS6s1uaGufBvoUQShm0i6/8w42FArJ4yoUvDtLc
RWvS03O/7y+zRMfrfQYzAKv8ymT4StAWGGT8kRRaH/fBplZ3pjVCNs9lvDPr2swE
pj6ji70ZIPSmlogYTbklvbu0DapESOpkFnkoJ5Ut5Cq1FHtu3Y0OM5+usYTCRM+4
PqUXC9n/Ax2AwhKL4bFCiF74Po/0xGA0MNTXf/d5jGhNiRJYPd1Dh/Vy8k7Axo59
s5i9WNn6qp9XBFGSnCftCHheUX5R6dCsVXdG+40ssid8WGXSZ/g+3pvD0pgsnn2/
a6rRw/wAqtfCIkT/StccI+rsvqWtJsl1qNUPXZUd3A4z6RXfPG4FrVORPLI+xy8m
/1RjIknW1IkLv5TNei/JjSxc4uzXLmx/iC04Bj0AO2OA1Fr7n05U6mxq4HDVyYXQ
XK24itYxmhirQAQsKtDMORrbxR+WTlPh5w9aj6Bmln4cGQwN7i74sWyfs+p+zxxJ
tvSJRvkyN+KZI+SoNHQvAcxQUP6/7xa6Hyv+0iEUWh5NxXG9WCexnYc5SbKehFJ+
r/YlnnmNYUtcRRJYmizKcMKMLEYL8zB7pzM0JRjiJnWihZWBMjSbQBMxWVbTnyub
JD23wu5j0CckGFmLWEEDjENgMvdBUm5CrjGVvYQ/fKRBFb0zRsfrOR14+2M/Zb2m
yObPa9cO3HQE3HFU1KP3T+3VkSXiD37SPlBkMtgGTgNifhNWA38L8vyG72rL4tuE
YmFWZKW2QgHXyr693Fs59oDiqAXS/xeI7nPiWrxg9XSOhEAeHILWGGz28XooLrQW
xlgt+xI4nisntQpSnVaVfk5Zl8/8NzpeWU9jU85SgoWWIkKYb4tmT2bEVNBV4Hel
eZG7DQwMYYJYtYRSwRQQnh1jAhKCwbrH/pqgoBp3yHO/HggnJ1iRe5UuHEeSLvji
x7YhA9lN6DHOcNKG4nEX/Wo7Zw7i5+23fGxL2VO1q6zk+z2a+KzMQLXGBXvvpHxU
4P9O65KxKM8snQL+pHi9bqoIUX9fPeUXd3F09pWW8RAv56I27ikptojoxercpMmD
kArRoNIXnuBNpFIi+BElGNVHP0erXnAiBNxyzuoN89i/rVgKZkr39YFeaGQO3aMd
CSuSJ0p6HJbBiEZXqyWKIqlVZeD95H7W1v9hVu2a/us6Mho30UcTE9V8Bb15EL5X
SSYuiMF8NUoRyFTUREYqRBx1DNF/Opy7gj7BmCv0t7oJC4ZYY3q2LV+UMQI0+fo0
vjJgFE62La+7ZH8YjgaXorXwyUFaS779JFEBYcYxBIfXLzZ01eIg5lHRHgTm8BCK
eQSKLrA26MVba8CImaVUM1C86ZRK+uIBOnI5iwZJsBw+Bm3PVWp0aDXzqTB0YO0f
eAovYaCLKrB2xUtR4zF8LGXCvSoGfPkEV4FQF8J2sN7ERcM3yk7lM0Vsl+qN3Sf0
JteGcaowVNpQqf7sCSb+mAVG9BigNfJamZVMUg5kjYCIs1Msy/V4t9StJjmYPSFz
muU9n+vNVOwjMxuArFBspkPABBhkobTHQWo2VZ6A7CvMzxJdBOSnZzslYOL6FdZD
10NrODxw8/iMTiz1WgBfkC7ikO2rsZYnkXprz6gh18iEtfWdizs1SnSLvbutbfCd
1MsOjN08WMwBXV8KhUheSu5pwkPfAmDVX+5uI0lm3re9jZfV0B+ooLlNYtvYpBT6
dQFOjvJKTnxdVyGyXIFPfbdTfx9wSVzO5+EcfV6vFWVky5XQcYlOdMfREyIMilKl
Rno89DXw6OqRnwFTyTWx/bHnfLNWNXUbc08w/XUJrKNxSdOFFCIdSChFQ0nGMVRo
s63i+a9cGyjMVLFA/FLal6amcwR9Ukw8hmIJRjTmIwqO0StNXuA55Zlco3J4CSEU
zsO86mPx+ISKhN1r/T18kTHtmRTOrekJWQ8txViFwB2Z/7FX8IDRpG//sbpoBfGm
5ne9ZGDG+cJWUf1B4glGD/bYQYQR2Aj0SlE9QXAMW/np88Nm3uz8gVnCxTC35D7K
rKxOc+NvBxat8DH6ngOvt6Uj5IrLFznP70WfKquxhKk2+dOQWreAWMGtr+XVMEil
GPpc2mV5SEzJFWlbF7jQG7vLhaw4hXmB4dYbDbpdodIM6i++0cniX5hZnMweXP/t
WwYlqze9vsoGgiouSM/Q2l8SPEkGARFo1x2Uh4aJbtu8EfVk6sz+oYVPVac2TmsC
prb4myxDlsBqEt4uJ8stutKFiE8G1pZ8VSfHNAqRlHAa6/LJTXqrXkr1UST32Xyf
ku/nr81WG14M97JjfuJlkSRTAKkRoz43OojHd48X8uoN1LUdTBc8Dx/yBZdBWXcK
sKgxNxchI8R//bbpIw1/50zvsz1Ob/EzpIzF4eGD5akZ9AwjU/lhx8ZhF3VjdBd2
VUxa7cnoAp0qsWsRpsBDAcblZHO6ILp4xQxZkOz+GDlFUIlrs9bR2AXkD0o75Z93
JcjNLpBguOWwrKT1So7hL4iyUhqBuvr2kRsHCxTkhPeXuGuLjsJ3wuxQNr5Jebr2
qy922J0lpNRilgNLHeEIzuHXMVbM9gAPuqiBn2SOCFhubtIxkwbnlMWEZtqppW3d
bFpUF71o4QAH+xfBRp7zjmi5zSqoVqJKiQExiW6kq7hlQwscBkeJxtHAnnvtyCSd
+u7hym7RGCOpQYYb5zi+sO/wNIjvnWrSy/p5/WWsBff4bmybG5HJ9nhX1Lkb2PJn
4+65bRmnsiJzT/F8uAZSFBNW0cMZ1uU9wNtywIn1vViZEn+4lJdukny3DG4KxzSj
C6dojrRbtyihW/gmeZO47uRCAVDEcJWWYIh9cMTCG8VgEGe4zKQQkSBmv2YpDdj6
It+LGI+dOqgFF7FdOBQxlecN4GXl5ALaiPmhIZOO0djnorxmbcVRs+7spopUqZWQ
z3Y6B83pPdfd8Cmcwe3OMg4hvmgsxuEY2mtA9J7zM9OOEjKWZBV+FM+Aayv5kGva
XbzIQpjoqivmyN8zChBL4tfoXQ8b5BJ9cOTMXcYcxjAw2rRcfpjaEjxFcCXfZkce
1piZsWlpm3CJEc7chnV6QaKC2+hXNBoWWQFZy5cb35eGjyQ1tk4K0VmPe3rVa06v
MJcs9fEzA5S6qwFn6+RbHbrZi8oGOr+ZP9Tof68C2LHG5XcYDVURPxDRGSQBbAZh
B5QshCBw9kd0ZYzMS6Ypb7WB2gCfh5qJLFE93Ha9kljGNc4KXxcwJQ0KckWNYDqn
LCPYklJ4OMG/nRD90e+AmglscfNDeZTCPy2wiEdl5Kf+KXj7qCoEbL56bAcdOOIe
Yq5f7q+2P41+TEgbpxxfQzhalVBHpLwz0ML96+5149DaYbfA+kKXBVWHUv9tpmV5
UQNPevQKZqG9NbQSeGAjkYYjH3e45ww3BSBeN5QVNNeVU94VIftXW0P8dCN6czcw
EmvNqJwAED1e5EA5b+JQ5QoWN+2fswCjrlzaF7H6+Ouzm+cpTb8/V753IFXx4VSw
jKXoKDT3Z/fQakeF1FpyFf+AqNLfLIoDU6Bp3PGhTDfi8649o1fkRwHoRFNL0yrr
jnyjvGAKHpkx6LIUSHj7xfXfFa2IAVCmyXWFlhJPyOP34QPPqb/DylB2vw9vtVDP
Ndhmcp40hSFD8bSrNWFZDN8jm+cYnk2P/vbdro1/WDx2sTH+hhus0+gg3Q3EZuDs
AgD3rIEYSh7VcABx6Wuzu866C8jYxVB+ade0E0vs4jln3VLt67OPTs+Sy+o3aOo9
Hzai2IvoCwXO+4pb6ZzijPrUJYNN15D8HW8BevvvcRYSnzTPMFvcmxmtq4P1MsdL
diL4L2u9p1ap9fFnGm6cb/HjAqaO5yWkRWzlHECokGDKY5OSQOjPrLJHUtuZFUXf
s6rYNQ/MgOGf2k8oicIZT7wC2VGTPSp/907lO6NKzqYbnjA+DnmoslwHh/HLKGO2
efXDvCzUwHMBD9wTw94KOmqYpGxnYQyLwoslCbwdwP8rrlIahKKa501mpzH0YaB+
KzmBlR9DXyup9k7LHd9j07Bf4DHvhMmDU/sIitMU4gDOaextO/WWa3f0fUCuhAp4
bg6Kvl8M2tAaOeIVpfRynNLYwMndw8n4n8aoQmuwf36Qj1lGH3sP+WdCop9f4rCi
kdUrXPbmELyGSIjeJfbXI+PPOetq07PqfZET2GODrJ+v4H39cuD7Pz55V75iRXRe
TQLKjvxBPPSyE4TVm2wSnxHxNcc8/qjW4Xt/PvezYuCpfkyElvGfZ//kPXhZ4DN5
GHWaE2r4ftmSeoCFJXKdxTISC7qJvANE80SLt+5NbdGdY9w0w6DMBPveFTXrGmce
gcJ8gkSFlwajVDpOQHUDOHlibG78hpctHKLx0jIzJrPnAaaqVEQpwuNXL2MI3fXN
B/C49xSBLDlUJMpWQCNwT3+fi7RI1+o2t9KqfqA+wTJdqRbDCgTFEKlIm0/oSKoL
7YOsnuX/W84xBBQ42H/RCZXffL4Os2QySOSZGpMXemL9+z8V/oNRwys9J+SwiQq1
CVYMOL1kJ6pIU2qAuii7FG5bO8vlfnoOxmiqhZdg5RKkTfumksOh2mdLADxl72Qx
850sRNNIqULFlw3NPVVfcqVQ0SKw1cJ03CqYEF5O/jjBufbP3xzwvbXmRyELVaJh
+ZJvwtNtCFeL4AU3eWq6Xd+B23HWastr+H+2dBDn6D6cvO7iAZF8FPqLkvytn+k+
kQcVmGflXuy6Hi2yp21ULJ7TrUMWSlgbH5NRwU91/bFkjb9WEhK5fCWlmuNbrmYS
y3U/CuLQULbZCWdbYp8Ymx8hHhHNIVXwX/TBQaN/DB6OKhMSAvEy68pCLFXKWhqJ
G13UMkN7gG995lUZfMCROTFoCGi6arxeDuAuZS+agBmzluJba8JSN5GJYiP563pg
vPB92Rzbi7+Hnm/eDb6qAZiRKLpvL6jxmYFuLCLOsGhKDI88eyu0bZzKGj9s+Rku
KKoAWPJue/2GZMpbO3a/DaW3GDhU+G4sgu0Zb1R8OSZrFSLxwn8MJcY2l3nQp8/F
0sxOkoJADhiElf6MVpRjlSx+awN3V9CjIYtWDINSQsrFSEh1HMXzT9+yGi6vQ2z0
SxyiPkt/LvDnHQtVZ0RK2KaPyVIJODN0hqnRkdlEeTXhs8EOkh/FuU0Z7KLlXt01
iftIlVqxrEFGgIGSQFg92/wXiLE6wBQUeXAw1MsmPkcdL2VXfBOVrQC4h6QnhTxi
VqTS/GWhhTMNe8Tt495nsPGQ6MwmnUrorl6bbHVreKTIBdBH0Jz6GXfulYYl9OQU
TAmeFmgY5FOIb8Xj5LZdwOn7NEDsfw5gdgqc/wdpiErffwDiuAc3Sdu2IC1kKHri
fVaP6zuGf4tJiQ2R/pHclpMATlEkC8sRSi180wKjMh9VcG7Q1iRJfxTfuVLbA4sR
33/vTrguTO3Zef1tJyOC4Fa0gXZeoddnqrRAgFGJ1/rfjY8IwihobbQQcU07TeRy
m4LXWLjGSO7cR56sXqPChUYES/LiDk3LyZAoZCEP191zbQcXQgmUzfrascdH8VI+
qg3DS+7gKJnXxo/qPltPAxXYomnMm0Owi7ELIa6BmIXBwOnzcff3MtVVgdb0DRMG
nkCLMJ2XpXVA7+F1XB583mKQw2MuXUPaznvqvkIGEtDcFwF2KDUNqi80tCIWBsrK
a6Dr9U9f63hsL4MpvmMFPBpKr0FlPaLGqvHwildbERa8Wsl2klT9WDDUsghsRNhF
FRhnptkJUENVXiIMC4scELZHdfZUQbaSceP7S59G5Yuyjk6pofILrYyPijuiO6nK
VaOKo/0+DC2kJPbPN/ydqRCjWUOD/Zurw2OWx90BgV801ckXn/lYtnhGGSPy2Sep
d+bsqoPfBrZXIXdAShHxid8Z+rRm1krPVgIIeVmzBO3heKDAfsCDHVqqfV4vPcrW
3Sgt93FuoJt7e9LjQXhYNYw1oDaDb0GasXETU7uEYJrEs30oc7GfUHGScfZios6A
H4xOvD5iBiO1T9wT7JbJP/brR88irWZnOtvqSZX+aVAnnTgEi91Ey8biKt1JNHCy
gdFIEOyePtzelHyiaQblQWJy4b3F1jTpUpLk6zSNueoUKGT4Yq1iyiMhwHqlpUx9
YJnZxONHms7TVJVxIb9CvvcuipevWbvbRu4FhwpHOCapUtmR0WI+SFIWCzCvdU9X
KfaoyaqhWAtaZfzqe4ZkHZ0zyM0ja5UlQvLisMpVYG3ynoxs2tDqoHV2SsFnrxvz
EFQ9wWxyN6DyiGnXdOOWepbUv9kqcKEXSO5wSed43138nhpidgp+ZtV2pJLnuwtN
ZJOrrX8Hs5NGPJyCHmc7xSXrSciYig4QO3igDKmhFM1xHuDMQ2htr3MuknOuYGa4
tqFjEEeoUfx2DTzEtvqVf5jqTCqC2JeO6RDr+y6gxME5T4sut3ImW3crFSdIGgFe
kaUK25MSiDEejz9c0ivf0efSRT0FiE+PGYGKsST0jFgCiK2JVUMXiPUdBIMw1qOX
T36gjcQwZjF3lilCpDc1XPVZtTHDpYkbq0vkz08RHb3JD8XXVeaZ7CQlF2Lzm5dy
n/AtBOvVb9dN8U6KsKy8uF9VewnfN2ydlFZoYu8CxROr2JzVNY17QpB1sk2Wh+BN
duILshTeVSHVU3OcxehWt+MxnPqOhhxBfSik6BnEnwEtvvaNoB7eSMGrj28t1V+6
+GJLBwQ0A4qmlA4xU62sHns9Axw3P9CucLMephS1gqd7EYeKFlW2lLGzss7CTTXh
TwW0oGbTW+p64tPY6aCxZNEfYhuAejzEZ/fHQ3uqyidHuZ9cpQ3cDIHRj7EVhCR9
rhVDAyFOxYIf3h327HxOXMQh22RKsqqHAvAA1IRWIdgclijSihQ0oTYabXUDNGyk
qadCzmbOGDDwsKkFxizdaKnhJYT/7/DXtI1GPe1fZnmQR9SC/lt4tTNkB5Gnw50P
59YLaYb7BjMtLVR430x1M757T2XUtiajvVd7s3Ey4zDfNOu1mZEcp+e9Vdyx4e2p
Q3aLKmkTGVgSbiFQGTtnXFUB1OYo7pShxEEaHFzeWOHRu79fkX2BLbEZ0BjIl7ON
BrVF0Yrunzlc6ulFx3OnYzy77yDQ4TOaf4LpYjin5IA0l4uBNTTtbly038KMa7Py
pxgO9X484wlO7MHlmiee1Qz8gGOHUS9goTs6V9mLfnw9Z/Nf2VznPwmfVlB9Tpcc
Z7st/jT9CsAVUbuNeO4rShJwa3d+7BUozvmcbI3L8N3i8TYfcF6PX+eZF83Gt2Z+
C9Z5Rd+FY8ioYgCjwEvMMSDdi/tymkvhmY8XHuBbJ186XyWJ1XEyoLnGbYOMVD5r
8ImUaDMYfY7LzJeX17OnePpA9/Qt3VL/kqSqHrlGd+uNTK9Grcb8ItTacNG12zfV
O4e9K9oSbLpvfPGpcSA5SLnoxdsJEQJJoDWMruuGxjYm+j5vEAWdXPuimi2Vi402
GxUYd0C5BIzX9xvowC6ZHkgKnRY/YeVE03LahLctEyddnlXe00AcEmG/QTjBqDBO
DeJBYR6zNOGGYjEZgBNliWVQN9rIznwKVOx91++LpAeTGvWIpHhFaZVoXEiXyWUD
WNrBNTJSmHEvnqkypebVKYx/t222Z32o1FPyg90uc9+fhq8bNPGujGZAaWm2slIQ
JHXYWpxRUrQSC2LMcIJ99bNQi2hhPxn/3tFG1cijW5vRoHvG1sU1A3tzhg2hjj2B
daIj7vpNzuWkvSjGmuZMopImNp+V5AN2Bix/nRQGllh+2LWmyBA0CprXB725tSfs
Tipvc7sawMC3wB/4HDxQAtJ1GuRst/KfwDuDVFb6Sc11Hl6CEJBmnsKF8V8E3BAE
f3jZ0/ulk8R5TCzUNefMIV5ATekM+yjVOmnu6GlcdAbJuaxfmxDXsjhK2FiIzNQr
hGddcQm2EZ1RXNytrCSLMyc8ziSeOCeVYtdRPnV+g3wXyR6LPFPIjEUo5/qxKB73
6NflHrz6my8au8MfCcHuPRvRIx7/4BeQPrmpQLeErp3NJ9e8p5GVZXtsjuPuilJ6
3UWM0jYJ/xssutt2xhTrIBhYnQdna087GEZRrAZAwaqUmyFozZ0l+4Fy5+fymWEH
jHWxQk3G9o8kPSeqgMLXziXzXwn5psYsPZXvOxTyqBPUJX9OguvVFgk5LvGLRsEn
MJ0/Zy9IjnZQJfCTY/EhV5v7kiU8uFuZKKPFPBFbrMWpVYLrWVDPDLDA9li/6uru
ozIaGSgCIYgh8Xecc7sR+hkX7aI3WJ5wJ+xSJ/gILffCIgvmwYcx2HDchMGCrIiH
3gluwRhw9p9aN7InRr2fWjMONDrLYzyIwVEVWtObDRIhDAr5rDfsJddqOBBhIxnj
6ZmTnqxViJv4J58owwS9ytseRu9e++M2rX1wX6MOo+YIpH3HTW0GvaBCYjDYIKOB
Twh0+A8YO95u1FfAIScidCCqhu/3Zvp0NPDFNS4YRbdALeZmYhsZv/7kulPHSxPU
Jw7uAx9oxOWC4eJlV6L7gwWe8wqu1ZsR2wM+CcQjx02Uq06/xqXPBotBPU0zgRqW
joPQ/zy+m5N/alzx1n2F/nVRSSS7PLStpcvCfVUzs7VmtANsUjJ+J+DlBgoXBAnQ
/GhD/DQU580zFRc+6Url5y+XnCbyYtqdLIg/8bT6XGSkti9arXY7385wPXl49Xs2
wUZj1cnj/K4pfmK4t92zdiIKXL90G6ZN7pyMsKdprd41jX6hygsAujwQw7X+L86f
TJAOL/jDT4cnmf0AYI5CVYTCOroXLnEEBGaowWm5C0jVixg2TMqZuJXPhGq6c4hf
eO9xLJBzXAv6hOc+WWJtsTGOXSE3ikeln6AHGyXN7zKnPvbP+4O+b6ho8Y0fdKGC
R4HViBw+5qH9dJvWS7tEEF58Q9Nop/HN9YlG2JvBei3t6ZhTzEsszWeSlXNAVKRA
Uyug9ifRg/sn5BKvmFWN4JG/LJQdIkeoSqoLZENJYfeFEgh6iQFAAshBfH2Fkr+p
WZJ64L8+dZ4vjSMpGYY6o4FRcJrNSXIpAf1zkeXfvl3OY9eKErs1is7IJ/Qj2ufD
2PqFp6CvIBEflPAzYQ7KDUbyh5x+/vm0yd2gfUPX4f7FLX1wISEKRvW2/Um71xUc
ClEdOvj3sDHjVa7m4SCQA5xPlgpRdX3SUURno/LDrb3S46xfCAEmB0VTzoNc1M0U
T31DTTW5n92L22Tja2PwvPgTtbaWkhlGWY7xTGfjG5ABzm/RPthNsnZcpzUohfAc
/4koPFrnp7BdVoxcQ++VJ6sUa9oWTN5N+bqbogOO+s/Q5W565TW+wq9d2zAll14N
2M0kmu+bnXMLhrnB9uxXom0f9Wvju7t8YRCGGC7Ex3cjyJ/TU+96SdMzK6Woue1n
av1ae95xsYrJfj6pns6WHOz57nOjZN5qAny+nEwO9CiWKmzOvI1WucLjt11B1BZ9
CaiIb7DkzxHy+5We5ATNNpbe+lQJVPB05RaGIvcG3XizyaXbChnFJ+N7Tygstg8j
aMCPeCUikNgH/YVkGfdsCj1Ez4uS6P6pGjMaTvMpJVuiiHEtIjthGZz3/mURdZV+
NvihBkG5i7ext+EEc7JIpOFkJpUaMG7klSdUe9MVHWIMedSlNnMuJt5VtJaRZtWQ
K3N2zWDJjxNDcwyt2DC5tRVMBa7E9OCUJAOlKeVYm7bRRehuxl3X/GZt8rhEuw9b
6HW8/k63pdGOSZ8V9aExCc8OKYavw/epS8EjLKjC9s4IH7jzj9x0R3ebsuQAHIAV
P7LFT5YfmTpAOXInN23C2IZC009lPx98B5kc5oeWa+uwV1d5FA8G+Jy+bFP2BOo4
QKm/LLuY4mtfv6sSTWgbvXzjXTheuO9IM+NWcl46Ynr5ZBNFuS7T49tD9cWwQQSs
P1HLxU7IR7LoH0mR57a1tvxt4W1cwcfgH1bbE1J2I1OlGqXMjcd/SUDrpyp1+0Ez
uJj2IJ6zfmMgv23hEtxxi0MEorSPMs/ld7Fzee5dT1RbVoOUcBFQEcTm+e2XehvN
PtcbzQrtU6GZ+7sacq+oRvgY/h25F9X0K4XnZNvcNTwCO0IoiYf+ZmxoivLINjEj
vsGkHCxIux++PyDvF0aUch+ysWN6b/jJjWyNe5oaiWWL4FCPVRLOXuOU+6vC1kbb
59I8MLYz0WN4AgBut2pOYf9ojItWonJ5kLoiytk8RgNLMpq5f8bJlbWVnGzDvqJQ
kseJembsl6d4O2GRRtf3bRltiimAE9C57ap03O0TdHo9kCV3jtYLjK5vbhZX6lfv
sQ8JKmJ4GRHF9gY99rU+qEK5TI0rDbWm9u6pTN7RuiJw7IaomeNNvc9xM1EOUrHm
OO/KLt/lhV81GaYKLsKCUQr8IULod6ay8Q4dKSM+zZDKRswaAflkazz0KdI0J1BO
4/mhrqIUzNoEe/pzNaVlAVIJr9sZh9fB2vPpQnnEnIG1COsgY9ighHkseRl81IYH
Jo2KlY6CkOZsZvr+5u0UY+6Jdf/CeXNNTLWV9Vkh/2Eru0rFQ4GwLou9qJXaxa+7
GGduBs8aywyZBQ5xAggZPb4yKXdgYnW3aKTLuV/oRIIDQGDqj7cMLBvqKF7DF2N8
lvTf3yKli/VYDTbIdnUUaI+sKaiWZtFvhF/v6tw4meTCXF0UOcXE5ZMJlZh6SDeK
dN4tdQfnEhbrRoXpGoZ15cAaJbzAZ+LANGMzWvwS8k1DrJ/JywXFvx/nef/T1IHK
+NBkbVNkPYqwP3SqHMu0yFrdxCiaZChzXiOM7jaWFfU7WK0G4dsuV6FA1Mu7qAoC
Dln2svPImS5GQfpjdexJYma3YWGZUmYdVWpbj4aIFQiYS6G/vdA6NRtjVa0hlg6b
dnkBeAu+fUfgSHpx3qrd57YQt9fMXF58/mgQvNK7RLBQUcJPZOp5xwZ2iehuRkCi
rDoLg5Wi7Nomjwg6FHsEBmhmXBzSDdbinX9RkTy5ooOPZENFgkX+LbJSdUHxh02o
2PNOBIy031KKY5hdyWGfSFAJDNYvRmkZ/0jv5/BfqKkahc1Oq8c32T21VY/ByaSi
/H6R65ryzf52XlmHCWBuzlZhEvGgTa5lyExfpDCx5xHlfRFoz1nNjCi8ri9V9hfo
z9osDvoM1kSRSxellTXzKnDS3Hjrx7a7bu+iFMUqti2yE2bzie7TXcI2DYbEg91m
xzhQWp/ZG9H4OFxXInaIh2ZdE5Rs2/48y8wJ3ynPGKGXpxfDKjqjyhnuLOsZrZJI
do0N0mo88dtmJb14k8M0dD/kX20ipEhFFYyYCrxjteu8GCF9UI4wdQoXpfnU9waB
KpX3Mae1IqUtERZUkqyE98taCjj22aPsR9AanR3mN3DZM4M1MJN1GzkAmbHAkVVR
0edbvKxsr2U0UEV4Aj8M6yoM/drufWjjs54NINFfRHwgDCoXniksqYlwZ1Wy0nnW
sIKRGPlegNFkJeenpjRc0C3G4G0jswkOJO15aHR3V/79I1exb5btqtvQ19Q3KD3W
uQsfYO3ysMRNWqHBU6cq4i9NE/Q8UaxHRQV8UFA6Z9oGoeW/0DFoerQwp12LqAAX
vgG/vG8GlcNnF2eM3d2ezbHV3AQCgNfQ8MLQCOwfAlyHrAAYzHoQ/Yk/xpEmrme7
ZRwnvhxeRbY/4Hy6A1pemi/jy+jgcYvQEvTLBRtzl8jABgSQDcslzadjfUTcNYeI
L9z8ybb10KOpj/5+elPu96L28wXuxS+yuKyuTr6lNgw0ZxZBy6wTK7yMbC2KPZVM
ReHGKEwhcDrYberjBrrIqYJKUL1oW2J1Wc1hBLb8CVnp58+e0fdPDqL0aYmbkrx+
fF9ODWiJFIDqKwh18zDxY72CVV+G+9rnZPEAjA7RYp5s4XTE1d8VUHU2IE4xJGlo
Wtnxx0dVjBB7EkrwF+H4BtjOpnjGk7yHsCavvdoDJkH/V2CE9Y+kyUITlyk5ip+A
OKRcRg5mrtdtln1gcinS9B6G/qP+tDoADljEW36dxeaF59JuWAZL1ELOoGp/vamo
dBa/iujqpGkpFrszBczu1YZY2oN/MjmKr65LrefEIGRgQDsPWkxmR9tD/U6m3mV6
He4wT317zFqBdzyZVLkmCnDQxJUpcj1F3QOrRqPRmK4jZ/kpTKCrMviwnGDDgBFw
GqbZTfQTDTj6MBZflcaY2MrfgMmsBYuO0HWkQeJ6RnelNEycjwVIUE/mxBCc8tPq
F/0fNHh+33GRor6wyN6fufUGA1Xlx2SgOeKFewpzTi59XVYu4T9A1FKd7xbEqGQV
ZaVEQCcPlRiqGdoV9Ng9wrn823CLqhFEHXH5ORvXsHOrCiTagx5XqSSfh+x/X0TD
Tv0Ap3Ma+8iebe50joInwoY5+8+AMHevtmXMsMeRKPb1swoIKQyPpOL69JmnDnWo
l5fO2M4XMoNznpf/kwHRSb7meNdddYVXYeO+mN8qPvycAoMFNWlJpmFIdbtImrIF
KNilS+PwP06RnOjh53P9vKkZOoXskwbaGFXbzgO4M0xfD3PaSGB7zQK1Su8Sry15
0C8AFR1OzdtZCujeKEX0dt+MYz/uBX+CfoDD151Pg30QHS5Ezm0QNCu/cNPGSYwu
v08lLQIU0Pw5p8ld9TTB2AJ2MyZhQY/RC8wTQFuX926Fl+UF+8CKbMJokDojv7ke
BJGeh6IF0CAehD219TtG5NM8PYWNYiXqPAgssFM62RpIFsZc63iQ9du3Jr6z7ChP
ZYyfWEeYU9/hpaVsQkt3BSMticoG4Y8aiVs2c+5Gjkfkro15Wlo2mXIsJqQZjB/+
cRAtsZeaJ3Q1BJTfOL0Dv/+hXhGHXl9nTky7G0MCBJ3wx7j3CbBe44v0M2cCKCIK
srP7iOxjL7O/e7dTMj15+PzKQOGNAPBZyEXK6xb/iZ7hcuGAghSTjpL5BdUtKkct
MXMN71EVn+SR3U/grcJL9VckHStapLaZnf/i3DOQQ9O3M7lQQwTdP499XF8h7Foj
/6EnTGy4le32kebecSOP97lB5xLrHbNXlxxHH6X+ubts+8RghxQkOrSP6QgF74cj
BjYp8apGN9O8oofZjNQfL+5tQHyk14Xh4fQjFbH9twUaOa78c99Zof45taOsLJYt
5/HmiyzyJETqMt4LTY8NjLHrH+125456Nooto7b6/OktYTXlMy32VLCmEobcu9wf
HQBBgqEw/vfNv9ERVofFOkHsiKJgw9lWtSpZv6CfTiWJk4WDZ5dWNOvYVSwFfWCP
7W7bD3k8lf1cgq5PfgTKopFTISCNkXum6pz3R2KBqzrm3T/vJNp4knsHaQjDt98V
hU5wIjOrbMm7GkGuH/2RdREAMETN6RSLUs3bThxnc46CJH2BzWRFvxhnpe+jelFN
leXAik/oXbKQbLXjW8Ei8wCUT95S+ofvR1xcoh31ajXmq7vTf+wQ3FU7q5XuTwfW
SzCREaUZRoNoX7g/ch9uCvJR2xj9MIqFn3ZSaBIhEXSkLyiwcsxN4TSOVNIHK61W
0cq2rjZt0TcU3nh0zpzIV3IYqB+YfZ0oxdZIdscbunJfoqNxe6gAoa1dK8yq9woY
i2fAOdZ7RUDqBtfBC0ei3jWuX5X7t2FXL9uhdSXUtEhM5yaLvI8O+6slR1zIlXBU
IUpZgO4HiDAhCWNcxCqvbCb0XHOqXhUjHNbJ0y/5QWPlKnetuRqGWcTRIpazYT3M
M2ajnId6ISGGYpif7jB9ThR55TZp2Arw4zy/7vqdiB/l/XKrO24Zz2H7vMI+qtko
0DWwLz10OomRk1paOA7nmO+iZ7ufr9EO1XFzEJ31A8m/8ZHNgZon8vP25+yFUBPl
JJm21o6q5FcQEfSph2+KRRcVWALHXtgKiIUk6PUXMWmr4N1Oe5MkZKS6OHEMI7PI
79P1P8A1LElCaUULzWzXRaXLTK5+EYwc8Z3jERtX5aE5Tb9hFx0zvRaw3cVIqfkF
K6y5qThcCkOlWBrpPmMapk3h+ZLPijOojIoso9/FUafqBjVJsU/3YuPIxIH7lkSW
d2Glcs2n5FishDu8+wsou0A33YWKEmh06dfzpp4IJRgmwAk4+0j7wzikAmog1Al1
0teOx93SUSwBu9osjwgjuxPtfS6sWwgYpzxAy7beVkwMe6bU+iqG7f3SL+wKleHx
3N7pOJrsv/4R3dLSxomfD8ath++YCnFErZUfX5CfDd7ejtWC/JFt3OdG2B1+CnD4
uDZ4T7YAVyLjfhtfd0wsYUxPG63exDwbL22iwiu5p9mfioqnrY9nVOSxWLAfp3A0
Vz+TNbJsZHh4vWCnWWFfJw/cmv/ZqNGGf6i9cGQL017nPoeELYXt1g1+c2Qsy4xn
y6J/OZjlWATFIrx0V7l8ohzX9yfydq6ukKhjL9S/PNWStgFrYzzCkGxXcam6NnVs
Kt7Ql9lXyIUJHQMFIVgXREunCmj315jpCPiGk4pzDnY3rKOJAcL5Gsz6wyYRgH+G
yVGEu33oCARLzUCPLxpO8zxx0xkPupDOjUlflEQdw0X7/su0AfWARZRNktzl8euP
EK8rgAChpafSTywMRewI/w97jBYCEKUp2h73ycHXkD7UKTrVawHRDs8HD5INeFzR
xxPSsoIOKKJwxwZ/yhq3q3rcAZOxSlNBMQ8oKERW0FhdNVyW64VA5N/5iERSk2Mp
zgBFoGX8CZZ1XpBLJnD9KdW2Pns4Q9MeUtkKYgr+TXKhUlSWL2zLGRO+vz393mbe
9abxlvCfRHhapWkvQ8HB5r5Par0e6lgqH1ddm4A58QHEoicF7H+e1Jf92PK1Fbk6
lhVD7b06S7tKKy3T9ScJdigi1Kb5L46r8pLaUz9qhAMaPOUXT9qKDFqjfMM93/qf
OE1um/4V8PzKC2yK2qZmxbYLJOp8RyY2I19gbJLH60R0mFjpDNAdjMwM/+oAgi1A
cY/kWFROLpGg+kOmZptT2UgJ/kSGzfxWSucCimO4MU6tjMLpM2iXndrd9d6nBR8n
TzylG1ANjkowiiMrO2oRc875dQFoIN6MZ2hRnMonhlvzeDFMH9777Ppv7lTlsmbG
xZR4xro0X2lPOoXMENYUeGyGw2FWd8tVRXiD96pg5J174OqKN9/mj0LKWTxKG5pJ
QC7R3X2NCv6oa2nvpJfuB2MUvFT/3WBC0hocc1JJWlg01THt7csRtEf1C4ql5Y4n
158DrPfO1nBupuF10fbqkVZJLjPBHL1anFywy8lX9CX6KGv82TJvzLV24zTUVVnw
VLbmKlfn8vz8FNgZa1S5bobFqN+QZaDgeSEFfGIogbOEdvZsyE6/4DaJz2VpnWCm
/apt6I6ju0irWwxmXuMaSVjO+o/dznZkVqPAwt2KiPpbSgkIxWWODs4Wwr8RSRe7
UkDxEyZ4hwTFfmJTSiaAgH0z5niTlIsq4Vb5zGs8BY0nVsDmP2zk0lMWSsQXd3lM
pP0D97QubdAc1tKnQHkN/OtepPwW3lPx87hvo7DuGddMpduKR1vvsZOXcoI8okXH
HzSem+AYGuhtUlwnJr+VfnfBFg2YvDpxlqxzBdP2su+E4JR+K6TZv75CwX2Gxn8S
fzvUdm5peKogBRpe+tLti5Kn+oxKVwt5F8M5Js2wMC4it+jQ72YHOCaIaGPHvy+f
HBC0zTNXqJdHORX+xeyUsJAzCORGOiF8MkhUIowKzdvf2yBqWsLfR02MjTGVuZVZ
z/s9RgcEYYNlQh3AHOzuYwll+SzKF1r4rJIn5yejDZsIh3x/vauNS+ctnq2hGdBQ
GNCMziNbhXILUt9JCnsf4D1Sd4HpMPxA4okOHhnT+ULhmXhVFC5CALC6jsFXp2n7
gZogjh9ZrOipl297OkhLWm335KJEVQa0a/g38LpWyNwyiQYdDqKhS3/vChrZEC6+
D+bmLoeW4ccUN5BRlS+whIW5VrlnOH2qU7ZBle32lyYuUTjiO0f4mZxs2X8xI1D7
iRawVjLdG502GRSnJEBNu3K54u+WglZlQO43glqJt/05tF9EgiXBgmonTzUTySPJ
Myvm0mYQyImwTYt9oVRqBDN7//50w6Fe3G01D7z/FBRHxztL9i5cbcdwVws8oyPX
8xiNaItCxL1+ooP2UqgpwcQ+BEXkChlF4IYpFIPFHm+8rb3jdNaxhRu9ErJka84s
G7Ap/N2Zz5cTuK5Nuymgh3RCdTLGpaad2DwN2ZqgWPH9KCV6IFYsmU5kamP/JDpn
SwJehqPRiH5YhjZXictdDllXze9gFgZFwAGDF7JN8L4YNcVizOrPbBuroAKB7P64
tIvL5erTSKSDpzPndYHMixZfsEtD/M5Z3QI0R1cjJwaWZc7yvJFd8JNNi8alVOTN
2OZ+26EO4hOLHdE2Ts/ue6J9N7fgNScbaIZ/SyT9NCUULunblZHqKw8Y0DFVlXP0
4yC97gmnzUeoKWj+O53uhLzDa6ZZZqvUBIo4udluQt/gxQzCPtxfC7/jESgGHuTI
KIQCuT2kIsmWxIoIDhTrG0iOawXYQYI4m67LndGAXRddAe05cx7fCtCoXHsvkJhC
rN/1Vdea6XuJ+/3xDzbLpLe3h4dYPpyjnCtRx0GL08N2JbHgdAM/aJv9EamhFk3j
M4RwHTzIrqy+hwFCN49Dp5FVr7y5Sw7OQ+1tYbsZ0I/qRzjVfskKSTwb4sU/MPA0
1LE4Y+kizpcWFQrqherXkVy6zx1HuGCCDSSQAeIb8gjwImjoAKRARXTKkxSZTg2R
g2tw2h3M+r7frtZ2dJIxnrEOwe5TQrwGlgziFSJIZ19es6EiBclE9q5dEoVsSTOX
sUZrtQlKwZ8ZrYWYbzsGg0GVM4Nf5vaMten5DgAtBBI6tigvwYT+RdzrYjOyvfdt
09YR5KsuY14lIATyk34PwrvxZ1nKIRqmpCH3es40qlmRVN+Fn6m2WJlUfNPSlt+s
KXRFemr+TqXfl/7zfNYSzK/Uk7YIh27uC268QuFtz2LTmgYxaMK60b/VTFzMVZZi
WrZdD/1MYvZJx/MMcrZEVKWaXl5oKTu/ye3FEMWfhMgAUusqNCzL6RNq04yR81xm
vaS2kBF+efkZs4BYiRQLhg2p4BGabdCNflXzxb2/jX3Mw6WTe92C0KSAbmzso7Ko
U7GKzXms80c01g1igkSm5spHT4FNJ+XhYaFs1ayNSCFHBuQFuYtF0wOLFaLHDOVS
eHQqcEsgUMW6idU3i+ol2gsXmyddxbzptxaN2g4cLG9I0PwiorxIridt6Bc2RuMJ
O3R59Et5j9wCihjRv9G8FY+5LZ9ik6IZOhuDCDn75mN5VWhEVRuJIJAa12hPl8xs
Nm0WjRxWdAfJMNRNlmQup5EhvBunQvF9x9Zu6gLHbqhPOWQfi1zNTS3xnOxZ+YWq
3LP3O1NZm0Fa9brcfTghvAGk11lcZLYrp38+fSNKfYe2l5DED1xQ+JIyHmsqzSpd
ns1OOdXOTziVcLtEX4dzz2QSepQ0iACLA1t4MNF61h/MpCwNObEWtZo8cA87WcKr
xImr54834VJpUpxc6J2qR1cxkzi5otso4zpqN02kxvS7W8I1ByecuzBvp1u0j0Kz
0CCffRkI0eRj92KmtlDktS1bnCjVnbQdaNejwmkDuzLJ/2XTyfnVCjhHBXEIxox7
VBdg6HApkXNDdNWN3q8dNgy+azoB7ed2oJTE6h3qm9H7Y4d3TVNcNoCF86/+7SAD
1e/X8DeGBUXeV6Tc/z1xHD0uBAm+e9e2yZLfoWtcNkBkl7rcoUT6Aj6qR8qHzH2M
iW9pDWp1eSEqraONa2tyQZXPwWu4s/UIYPcDhNHx5ccLMmadYpHS1Yp9SsAWcUoa
Dg5cZaUo4oMYk8PnMcxumQlXSNGPRGFU9JpYqbblMF3IhqJNH0nUMCqzftDdPNZU
BHokdxvYu2HvYVMwTcjYUV5DPFlT28j5KJFH51hg2f9gTR6gXyJvpyGKkT5FqR6v
fGQ67Ys3n8C3fi8H197EWT+MMPS3jj4AxjdMUxOTObwS18BrHPUlkTVVeFmZQb96
KYUTN+7H9o3u6+jRqBXQ+dSKxnyYgmCsD8hW3UPPr8RLPnMg/zx+ZrlvYBnsIwZU
xT4BOVxk3CH93a5MISjEPVPwhCiareWoBlTYLO3dWaZti/K0LZiu2yjUqjRJvUcl
Hb8jgHCAXeviutlIJVmEeHzBnG17QvMzlz50HMLqVCptk8MD8SGuIGRqnSw8XY/t
oqImVAwRJuYkklpOGwoqPjqTS9D7Lxo6mBLykgOjz3/YkgIwXPYFKrAjtGwtgZgI
Wxd2I0ssvwJCWAX3i714KcW7HP/K8+RYooMTm6MJVj7WXISJHcH0yWrrzBB9w12v
2E/ouSYj98TAabnHfPQIz65i/quu2/0fBIwUy6UwFJBnXCc0T9BnGZQb4MSFt+ZI
YvDs5D9rUOJYMDLGkiX0oYt1z9LmjpGNhMESlqGx34rkcZgQtid8QqyKSJRQIh2o
96UoBHb9c6+WpNTzUGJKLJOZ/8VVHQWfBHaKsGbCn8ah+9I12TexiN3NbBfkS7lv
B3x2zA73asop+uDa8tKKKhcpQfhPhRluGUa750YGu3mHgpCCgpmtZgJG/Iys7Qmv
Op3SXyHUDK2su58H1P2gEj3wWu6E5KF2g6BZOPS7D9fy5QU262qu3CM6QqBNM6zM
A61vHOCPsUc1Y1sVEuG7dtU6Jqf6MD0UV5ICjMeNZN3udR7+aIqPDBSEaUiuFVXS
9RKvk426j/joGWD1YbCTf5/4djU+bgGGmoAsK4ZF5GRNjziq5xx7DJg093adLiGC
HmmYkEl8B5D7BbVqA2TSLlyurV1MwmfKZV57U/YHP2GW5EsB+5+1sqmiDhROnN9o
WuXK/wuN2vsh513dOnyJ7yYOPK1zRK/DTtd24LsUi8K4ZP26tgXa2IXULz4itsca
H0bAKRkB5uzArSG8/6h49nulyIaenALOI3r1zVzIyem+kg0YiWmZCKz2cIIW7n4/
K+zbrtM8vxLEMkmb0dycTuq2ramOn8QbACADq4VTA4/gcqRVZN6eX7PYfB/PBwhF
UWSHdT1ni86PfMrbC4SUSW1ikQsvXAovL/g3jcqSFVlg2KTQ+ePN3jwns2gTIkKE
kzpM8Az4Aj7/wUOnUMy1W8HxPODClhK1UGn0Xfr7B8QLP2ty/LnFBHkGJCXih5Vb
xynMqx9byYcYKnqaCyUws5jqdb4h+90r4hHSqoV6adKQl1bicJy1uWIiHy1CsOmh
4zKK39oPIpzOtT9RpQXPUrK5Rxq/fY7qyhPpNoy3sAgP1dUOrBVY9ISjrSkTDhvA
JR5Hau2NdmLdvPEPHOwxHAwSQmAkQtjyIyQ5XZIuZYqtiqabbgeqRLIofSdB4JGK
crh/K6/j+hNA3i1yoEo7JXpgm6QL9c6r0mSTGgD0iuMnimmEZFa/vGNWCpUrlda0
mUhfX0v2A1W2t5xO4DIRwuAG58SBJR4sv8sbtx3T/TTKIahdlMxuoFPEpXQjUy3o
r3Ovd9z/+p7csYRhwv4f/kN0tRVtAsO6DnVYB60egSmRjtcs3F2YaZt7bE0x7ktu
F+AkKDpkfnwTNKdHdBxbK5E3YnheXt/IO/KMpLLtmvMIGwqyhcTxwxLO5ZMu672a
tmuuE7rkN8ye03voZWBVINyLvvwEOMJPalbLIA78qhzZOaPnjyJn5fR7UKQ4jeZi
2R5Qfh+nbDmeKEBrTOkhjUWrMJenlVEf+5+peDctppk57bF03ZsuunQdlHxCWwi7
TjODxMcb2D1HDqHzfB+1PME76St/3WfsYcdUl0DjSsrJzhbJkJyqnHd+X93CPdr3
U3K07QOLlcokzQh3mUYO9SF0dI1n8EmYG5yXpNCplKu7LJikBu7+zOTJDG5UebRS
A2bVuxyCyh3Rhw1p17tnaacGkuzuNNxO+nvaj+osnFTsRufC5GiysEOFQnH+Y0Sl
yk+uNVxc1GXUC4jfbH/mE+YDP9TcyiIHU/kGjUsKV8mC+E95ZXdMn5uxswOfQTxA
kL7lm81gcnSIYpymPTePl9HgSgmOeReIODIWj4e3knTgEZEgrm6qB8Y1ifiF+CEL
SSLCse9+/vjk4f+s3ySqUGrTNojAAY2C+XwGSmhWrlJQA5HKASB+XD63CumYlJhl
Xl2k8ehyS7z0ZPptxEsDQ9Sz50rIkcjsQA5U/JO67/DoQfge+ow0lK3lS1uUcejN
bEB9XIp99VmQ/xkmEJhe7nmVW7nmjHr53YQvMaXA+KHx6ErDP36P8nR7d4q5xkmC
u7BpznRd9wj9TaxqstD3cnHoGb8ZNyS76M3vkFxE4iXiRwmSHbYKyTw1jrTLn6gE
oDZX4s5S7lFCsTze8ZaaxZ31bQNyUm25qiKLIBjCa5C4XNefwGyotq/wvZ3eovgu
vd31unulEIj9mvdCyt5bRs94JFav/AID9C4VEIj9So7nkYyxaPyS5FmV5WMO0k1A
h38LF6uC9tiRXUsXoytETmtm0BwbcEmr9vI7oneKrue0bNoLDxP3Oi3wJkP5FR2i
lin2/Ig5AN9jjbiC6nM91iu0u6OWhUUBZr4+jh/Tpe3847QwwpNeyuxn00wDDXi4
onsBvxWRknkGItDPnvy2bsYFMMxMChTv5XpZTJUJsUzTpW6cT8AgfDQO1L8RgPyU
1ZKJPd+vCqL2/oGJivYgSzq7XHXGRDZNONaF97V+XRuzj+NfQ5k3p4g34Qny5OxX
wPSy7CPGkis6KtYex5YGT/IwBsyHDk1Povmh7pcZEyuhqX5kjajgbNu3GlkWRIOF
YOj4QjfheIWoo4+p58Nv0uHMmA/SRnoXrQr3D28NfJ9MleM1RJGSeave1sqByfwk
v4YfPXusNlVKSTQa7lhqTsRmZEJcyEv6wCUQNgKCS5YSKDdQZz0iswcDlRfPSaQP
ZixbgM9njhwHL1UPnJNuWrlCTQlMqwQfd923a93RAF4oNFc+c6BKPQ+hLiHIbuM2
YQBBPdyjuKmVONiQ6FVDe2kX3eqP3PdLXvcp6C4AI/viPClBkRv2fxUEyXoqdziG
BRUfwxnS2FenYj4z0WFFUtPpHzxFFPOoO/+KmG/xZMSf0iIpRcdadJXLGSNDhWKq
enDOghQ13flOuOkVygzdaQjx5JVXkSAnwGSqxpsUDUWAXokBehAwWXpTd5twZL9f
ViThfEvsFwkZKQ5pCpKLPN194VJKnRqw5bc1VdBo4BQ/KCxG+WMG81gIfVUUe4PV
sJjU+FsaDzJClS8Zd4/Ik25Ag4XnI7d7MqddE7rVd5eZmbCWvxVzG/H8+0qyVD/o
X59uuUw04xM1RJ+JTG5tD3DvidJOmsd8hoRX2va76Ya559whJmL16mWP1w65tMKK
4CSPaJecWtwYhraIHkKrk6gGjWQmR2n/55QbM4i7NtHVaCSGokhsks5m9xq11fKo
3Iu70k34VMl0Je9CGfxXGopyS0esFkrK2OhWeUliGsnrR2OnCaBHUd7JTcuPg1Fr
Cp+4mmXYTtaZHGyIRQuV3CbMSRG4MyoorZvStEgmQOrzAYGxaqlWacmsFbadB1iK
hd9Lh7QQvHfl08YvxCZaVkPlk6pk5x7BXXsAcRwbOE05BsyOA321Wvgz5SR40od9
x+A/gb09C0mBOewYr+iZJmKODrV70yatuIgmzCMHmvnxL/+ui1bC/t6Pluoh1Qya
M6O2Dy+ZNFT6LNVIHfqj2t1UQDjQqePqw3Pc75vzKovJmjieAzDp0/KVxnex2cwg
TgBq/xGbIFZnUBOedJ+gJWEojRxqivTUNFGke+hR6F7ZyEhqV/wPdls/cdsP8mlI
YHMH3M5lEzTYqbG6Cjv+uahjw0+gsCMBg7FH50kOXdXzCtJ9cQpHHUUwEZVAarn/
0vsHhV6mCho6HNDMcid8QvH1GSfIxCeEDQQtDAR20V5M5L69uTqhkyEj3yfhtR0Q
2NaW95bI1UNe96o5D0yfb56PoTEdlxv2vmldMFd8GsD6LVBeCwf26PRxpjZQaYdw
P87sRGN2YwaXKiY7EHbc+jhimkL2thvQrttLA72BMUHpucN8q7VNvTiOV4JDyrEY
CkxRnt/Q+W/ZR+Wm+3lQDbles4aPKRs0hDVSWYxh5nkm6QohBrkk1LC8qa3Mvojc
aKTTzciq333PM7uELcOyhqVls4nloS+T6/ZBbprhiehr6x/i2G1Wrtr+wtz4g94l
hTISuQQ5DFNOzxUOjJ46kbbnehd3j7+R4hZ96BVBPiouhnQ3oc5FMwOrXTgMQteD
GhUSkLUxG9MsdwXwoy5Ua0c4lMCjOo/GBlMPFS4MF4iQexB5+GnACDY/nYvnScxz
3t3mnIYON6l1zO9g1rI+FSdN8J3HrekUTepBolEjoI34QbY24b9b5RG5s53JC5XR
1DgWM0610fiiB4/bomf3oEv0QeysiEBQdX3rAw+QjQ5klTcCAVhZbsV+ekU5hMvn
BelwmEVcMgEJ2vm2YzIeBzi8Oc54lcYmp2C8oUavRUin7VPNaspVug8GH0U5NJvh
i9xYZM+Cb+hI/ScIqFM6q1gU9pZuvFDK35M0ZVrexratlGl81jZAFqaejvGVvN7L
8MiCzcx21ns00wyNrCdH5iMAZhtAr/4GqOT6ASvKZc1eu/Mw5dGG0pBdGBjPdag+
cEeRQp06/FqUPSzZ/My9eQVHZ8kpf5EMWXOeCGj15ZoByeCn2UN5/mL+2L6L+M0w
0R0V0Kw+X6PI+mtjlTpvcEk85WYUY//a09RADN1EEMLYwoqAJ2wOTXn7OaOIrWCz
oNYsbp1BFACd+MBPbysD7fRxw8UgapE1xfddGFdNxZVo/UNhoodL4kXxasgRO8FQ
Y338LzArFay+Abkrkd+sW1qW8RdF8fhvs1EQvf5+0vUREL6W1kgylNyt5FlCuODe
crXW6EFl+PU2zxeV2xuqvKsVSvTmUIWFXdE3umO1lEhCV7ovcOXK02jJq09lCol+
XezXOBw3VaTJVIx5zkJSzz2cmKnJdI6FNytArlw9f6XWSwyU/NqpdEePghz9nnTo
FBxbA685DggOJFztytylpe/0IMqbIE4GM76gLnWBEPqo5T1/klYQWa5gm+lPNbYY
1GT8EPfWg7FUyyHgPa6tYstAa92/8Lm66NQMCNKOBZQR9aL6mOkK6Xvh4x0txdtQ
mUnK/+WazkCliTB0vi/JSy+7JONJwG5/o37zdH7mUnuvQc4S7ToGS7F9ilF4M48f
p4t5phHtGhCvTQXrdOo0v+y4yheDKBLz/DPo31FEiKFm35BuBv1jYxYV/BbDLviw
rBNNOOysv/mTTvXot9l2WM3VVNXKP4JZI5dfsCuY/ihsu2lHsTT0YNEj+7ea5IxN
B70Cnok4r2X8XR29erU5eZiW7ruRjQQYX/gp6ZPzfA6tZ/v6qy6QigY22I0QszdJ
1gLmwtgneQvZ6aJNfKth7gQaXraVSJusq3KSWLqy44DtGbOJAFoiha3e9feslRlB
OU+DJLQMu0dZ9KxRIuTlvD9F/BNhVKfLnY9OgAv4LeNKWLbHfdAnKeIJt06IMMJU
IAB0tn1dtlhgAzlOVzraCX0qVoWDCPV3uGlYEKOMGrihJtg4aGASMJyUX1AKHiVh
gCNX2nuQUIYoek56kId3oDXukoVHCgNz9umW2NAtr2dNhcOEkMV+wc4z+lzNfnLV
i59J+gZ1SjEDledb/N9zUmFVohXiGmopIqhFqd9EWZd+m1btDUD3miZ7+eYitczS
TfuY4zdDRY0dBF539yn1HTb32g4DKAOfjFDI9YiobwaFNNyONfUG1jEAro4Mv58V
JsW3wZLeYTE5kG9TPJn91STeiQGXQ6H6OqApQG1QYCHRGkum/bRAO6gRrq/KvU3x
JtYvJFZqZYycGntIWZTu6Qqeil+oRj+d8ORUaskJQ1edcmLxp2lfj8KW6g6Zu6xa
OIzfDdvnryTz4cXWRLjPwq1aBCz9Woys1/2H1DMDTCQcecRVSHRAUfqVPBOA0gdw
30hIULuzJGKZBpI05Eo5zQF05Xg+hOHcEqtmGgZIdt6UW6318koA4bNRvuFhA5nM
hTZGknchPO2C4VNDQKjZi44wVarDm/tZ1OnmAeV+HgwLh+8jx+PbiXCUdUbklQEC
IT7uQrnpd6ZNmEIlb3Jw7RjbDZomKf5cbV4LS9DJZ9Bc/63sVopb+rNMay0CHuXj
WIuDDHPh8Tj8Qt2UhyISFztZewt1QBdBhiq9G/Tpllcw+RJHnon3xG1Pgtsxu1Qr
WQzuwqoP9zKTiv6G/wEFpfA8ZtyJjW2wd99b6IfFgAElO2XNNnt+LkgOVzxmbs+S
atFYVZI6998yPC3hkD0uauy6IbXajotA/mCj4rQIkDEeOUJ3x1oIdA382Bz/rwX+
Ljko8rmh6XI6fKH3yHszgpKDexdximbWQADUcdKMTkK5bKjTBwmkzvT9HPq6wNBr
8kVfUdv9xR5rHT01k4DiafVuIM6W+tbsF8KMdAmKAyMT62p+yM8D2do45NACF7Qg
72i/Nx5uOj29E5wvylD6FF3jRyD8II/rjzDojbfw2C9eFw6MUJIXv4UA4JFgbFg/
gGkjnc4bs28TvmfFDnShFOvIE56v+hpHcgoWlRRLGoXJynz5qEg0cRGt+qaoti8W
rPaSMAey5qjJ4ApRbOBKTrur0LVmCJRIQLhRZ6jq6qRneZMZ1K69bLms2BzIrTv/
Q14gU+mtuMyrr5MV2agTeJQVZizvNwJBBy9nA4xFcuxejVLgKjdMdb6eXtbQVf5H
Ybko81fGC0MWExZAdaGqfUTO/3rEQBxDPwdIIiFpaIapEyBUy/dVpf/NwZLNtVoW
ymAX5OSseqlrFg5dnAXqNMwwUNHJyu6kJ1sNUtxqzG9rMoIx0DBnJ1ylQdqdw/1Y
XMRqW8cBTLlIClj6/nUSfIT3BYS/1Cu1zYU2/0lugwZmoN7zrpEVFxhXg7Nu08Bi
XJFbyOZvahHLVXLdxA2vw4hVzDxFZFNzWuG3Wvwf+1DLwtxAuf5cnYZJai9utK9g
8l1yLv5812DoWQOF7+KjlerHLI0DJkw2UWwbVusivHgo52tsYFtu2OcVv3SpLjAg
ip3f5Rs0r3Z3x4BlH7hZqd22EOBI1MffBbXxVAYVbzHoFJwAAM1rro+MIpMb+P28
6JJwmZS2JE0K36POWvftG9rmEpBFYrGRiANi66Whjpmu3By+FxCEyS4b3NIqeaY3
Ty6P/Bx3qRA3IynLpkBORN18IYy+yvJLdBPVY8ZMkdgrGDU4QTMYvUzoF1flpvSY
5Yo2oTdN0yP/iR8cfN24KnAKTzfgR83V0U3qkt9q8Z5BB+QH8c/Emxdg47aRkWwX
HghiPh8jzReJxGSnwM1qu5YPtRm4ENwH47U2nRLmvD2x082HkSvuwWBzapdWeBQj
XdY1ugbNzuWtZ11TB4UJBT/7bWGEPdOLHsssJPW+BP1RAmEwZIecH5LkanBTCQDq
QryQsnaIFjWaew8iijCmga5v3VnQMZoNjAz+5m6Mil5vkajJiWsVVlQv9oVtwt6v
bBQtTCdxlLugETTe3PIrti2fEpWTqsy7ezNYPZMRccrpkIj53Eu0cTqBVxgzNogg
PZ1Y4dE12pGQiLB7pJVlEJK5JWmkRbF3Gvm7+WO/hJQL6071fIlPd6M/2ELqeY0/
zLk9zLOFoknmkHTMWb2lKw4ZUJ1QJlRW2+dAJ6c1HL1EegQkhqSWmb9eGGA+7tjT
+Wdy8rB2jHTVkEhblTNo/pEdSxjnT6s4cJ+cFvRAtbbA6XRGr3JeKIM94NsRlgdQ
Lcx8iujfzHz2iXaNd9/u4ZjGTNPB8r6MSWi+3TugXAoVvdJrTDiCr2RBmGpMTC8/
TOT9nGCCW1fnGW1kwkq/e+foJXd/A2sZ461wt+0ujzSPuh8Yh6AQO0Kwx6JuE6sh
GbFSurxU0e2Y/5cWI6uAZQGhi3ukU6d7tfa2rEZSXy9Isk5b/MmCEYQaytvI2X+r
0tyEu1I3lLDxs3Ih0L1hM3bc7W0ajl6P0H1RctJL8VvQgEHCLZvDIL7lX/2cHiUg
90fn4/muI0X3UKWEtkUHKANl1YlQB39dwhfwrxR81UNNNHttVy+eyhSBW79hBzit
YQiZU3StdGU3O2dx22N0E3sNd9yzX7cRfOemf41xgEI7oxfWShjRsbPEzQIYKTRX
D2woVZXDxhpq2tBBn+DQ8h9kX6GYz0JnwAIDQ4O3VBzJftFRkyMJjFXlour3PYlR
pD6SeFD49qjW4m1Yk98X6+fCWaWq66r4/nPflddZ/WkLwr4TvX/rL1ci4eI5kBEA
3gCouDJdH6sPtFGHjyGTYckUHqTW5rGhqQhWnkonIt4K99tcKKDEifzlzKzEe2g1
dpgcOy/Bn4e3OG8awy5pztIJ3CCc+4r399UF3z4/7NpJ2+lfJNSgS6bI16Vjo96g
8EImYneY6zwDLUyLG1unoXOYJrX2SATezYMlPQnpHHnAEnYUFYGH6W0VLziY8jpb
bAGLMG7BVg1VzzfwpaGxxHOoAyQEXErJqNbOuFGOjr0o0+h6hDEYo39x6Zmb6Lx+
eNU3s8L8gR4LJqxTpmEMVXOt4Ti5nh5PnSJ8Nw4Hpgz8N0V0I1ycCkZjSdaBYP3J
AJ4zu9ZqjHh8AYA/v9gc+Ny7LrMMP6jZfqRnzZNme6gIBA5FRPgiiLUmiB4nMBE0
bMh6m8Dr3Cl5ohaLclm+En5JcK2Ir8tNKFq5rOjLRbDNb+xOo7JwAnvbzMPpDCRW
tRoTrLQpkBW0RdCKDINGMBy6wQ9XKsLVnTRvZsq/js/cJo6Wo1lXb5ay/andEsT9
Cs46wg2qfbI8rTAwnFhxAwUdRH1BJKXjXT79AdUIDDHecN/xyMIZrrumVlxYvXKC
3+6KcY95QUfbkWbPM0sPuTIrIR4Iiget2Ex7Fjfth4Mahhjyop7NlEkp3klTPqHF
DUqsq1X6MrGWz99Gai7eWcYbY/imCnYvNgRJahgvrO1FYsMBfLrTiF4rRps6f512
oNY0sISXDldrIPd7awEPmZ4B3WsYQ9uREghzoXethC8cyQUiOnqL3b+6qFU6Pfas
NdjSTvewHDSR/MxUyTULVEi4Z2L+nnFTvcxdxpwDwbj6kC1DzHtBcdpVTN+hTkwU
p+X7IR5LrGpPSkSsXVsPJ8uUWQTiCiSoc2NAOv2bokTphuZrTHRdqpWiV8X0tNDl
GNA8dEon/ee2KGNIG9RBfyWPD8smMn+M4QsO0DUVa5leWNe340szCg3U7DKcEIPY
RJs6jVjmoLZvlR6BzOAfbK9/OTJv2jU18ruYF/7WzkJ6fK42+hM9yRORXOo50oEk
uF0bcofoRLFTrodsP9qbThalx5tB+qzXMhSx+Y0WKHdO1KczHaqFzYulhOd/pCUb
IQMM+IK+OG2mWbU/ZK2f80XlQ1EC1LOQPMfcgXOl6LGKqWyjxGbCb7t9fQZ/0LxX
VnMIMyBN6asPPhF/kMb8T9pkS03VcwKx1cgtyqMe3MLSkMxOt9jpZQ7I6sXySPx+
FYH2YPbr5b41f0hDtFSvuiLJA6ce+a3DhZCbG3EOrucYx1pDNd/kkBQwDK5j/SFJ
EtxlMFCXmleCMgd9+lRVyWje9rcPG/iHaCceGF4y60dTnkcU6bX5XnQBaOnVt0c1
2alinIRTGFAMrklWL7NffDBrCq2VcgSA7Rrz7br0l2LcG1lvMtOzM7Yt8jKECM8w
Hq0GCaAl/YunmBkFC4JDzo2Gi/DbkIb3pi0+gILj1FGRqQdftRD+MyBO0hmYAfOh
Blk63wZmouXbE0GCUrfLTNk+veSQ9Ug9JefyQ/XJfDCASQlXrv86yolRcufO2Vmz
NUjzbakPT+Ao9AvWlhIb3rVYWRVcUe3tjB6APQscAMcUE1qWgqgk5PyKRCYFDJug
K8H5HjkQi2d1RqUIBXa4jgUq3/BCjR/W0pgv5lV8nh+I+GRdMweTnnnhtlqrBeR9
VkXW87e+6EtbkqrmBwjuBTQFLKzUs3iHhA6/ZHUPMhp19ACtBR5bBHzVqTJQ+Wyq
laR4BqtM8fOwSMN9gaostHQV40KoixMa0busyD89X5xD0ct46difZRLiyBLSRc8M
X02G3OKw8NazYHb24idSgmSszUvl4Cm99fu/noVKFB19dWnGgV77M0CbJtiJjw71
vgF3xh0YPxQpsdPbaO0yXNS0cCj0JvwP3WJH80xRlCaIBBaIpX46AFl2ra802Bxe
zD5mVBlOYtgJUrAvtf6WZidK8BQ9g+pqmPQSuObUuiKEEv4fz9xZ7znidApzmOPU
eLahKUTmvMhlErraCjD1xfa1zRappi8S1IpWfMsO8P5oCUKZj/XfhLi2M4d9xQg0
1BnRwE3K71sTv3VR2/CO4qRSGCCVQJ/+rw9icnTAQq/uBl1OZIgWr77MM7WuFXnk
a96di6USdCc667X/+bRQM7yZxiP70e1kNljPLqtoJo694IsAH2ammndsNxlVD9KX
YCztOtXAKdcCu4psrI34ep90IlxtqxktYrAakdXAZhy8Pfzniev7aCNvfbZne9E3
7khZXBH0Q5dyH6RzIa6MNVDyh27m6iaMhPfOBaxw0D36wvxgk3UNC1kOQbhazDGO
6XBlLQAfpEGONxDdRd0LDWc0MX3RIjHKGewtjGegrlBooHLG3+2UNVDqbBpU3XCu
3tOpXwnXJ2GV3hlAfnxcBmTgK2PnYZIcHWMgLWcUXVoai6OnRxDu5IkrH7p14D0+
JPpEgnwt+jrdLN9IXYJn6N7gd1pvh8fzqywB869VieXeGsvRoOonomZj75D4+TXo
IoKIsC+rzPtegQ1RzkbaS440vYnZN2sJRQjbnwPSAsUfEKTujdA/W4kSBhgxM0qc
/4UaEOLxhRZZ/baFMpEBuOFskc1EhPMGCqG+uPKugBNp0eKM5662/GujURAZR7ex
Cddj3MXd0nioYPdTtK6c57XPrCyAABiiTyIVACN4dLwbufwsA8E3q2mEvTUN8bFC
ENe0Axz77pU3mPXjpw/n93sFIfCbDyzDrX+1aGhN6xTndgCyXCyomKrRfYoibtD5
Q4NvT9PNjHW9kB/yfXIz1p4yX9N9w+PV04NHQICAWF38GFFNUiOMcFh1vTsKmPnX
brYtewiFJlHUhzKPTe8o5n2p2T1HSDRKLGJC8+aeAJF3QpJwNo+oLejvUB59qKHH
kId2paPQxQOo/h2OrZSgVM1fVDa9h7yPc6ghJqQ7XN3xrmzySLT3jdh7N1W/Mi3e
OhbHIRK+z4ITfWyAsinIa4NaIbvGdZKNymXqJZzBtLSI52dObAZWJFmznZltrnPU
KYDnQQ7Y9npdxAViyT8AWZ9OORlgGILY5HyfXeGeILph7WhbvpRmTYDCiAn3YFJR
3UIIDA6A+krKjl8pvqdAnq5itPXie18BLzgVyLwLTKu8JWXPiXd8T7KsXg9a6G5W
mRRsdx/YPZHH+Lfnxhqw7enJeBkHbY9zVykwYXPqwLLFZzVdasx9/NB6TR54GqIf
83Tfw4DLKZ/KhTxj8MscQqHumxvOe0EmYLrx2Yxa7dGDHFv9/G1wZ94O61Wxm0jL
wT1Sc702iqP5Wgqm1wHLEF3E9bpldAD1FbaHznM9GW9oY/M2pa9lf3wgTHazPJdZ
a+DfmSVn5cxcgEv9kYW35YTRC0Qq88ZiiO1TmmTJ1MCMKYlc6/zmC7d1duvJSwhb
VfuNz63f1Xs0u3m459wBOGS0Xq0MZTkXaC4sGmPANqfkSe0GhtP1Eq3c+tG74gwO
q754iDW5yR62V0XwRRgtnrNenTucf7/INguAXhVFXW5Q+Zo6VRc8wJxHmzsJm5ji
am7L1ANcoGKptsp/YTDypibQli4CcovxEXplj46Wf2xS01/P1bsq44xDHAuqevCg
2zjhOEaFRPwDRvjnvQV7jOM8lVbt/e1GQuLg3pyLtXBNoj88M41DekIhvAv3D5lg
uxfx/GWJnUYlNIbGb1gAWZClzsAZxclX20gQ7GPaGA7zULxgTfEtjeXWB2SgcLX7
cOK/PakMIC94HTDgtP/jFgPt2YLQalitC23hrx4OiSPVfFiWsmxclc4JEd3JdeYC
CI5qGD6I53YpHiYppHL3d6jlCvTKTrDmfQFZmEHEwgZgivHDYhfdI5Zx+XzDnEoJ
mcHxv0FmGz+A95TnH0JCKODGc+tywZA53qzE5UvM/56edOMWBqnZxTfSdWB5uHDu
cmsHpT7KetNlQDT/Kixqp7ZetAJ4+Tk2y2G6RyLidZ7b28vtnM7oS5LngU5QA5It
LoQKPd0U2PlS+gWVzyjo33A8xBpeIf6aVVcjRRWJaK1wkFmKjhIg11SLYs+RHaV6
yd/8oYJv3qsEIlf7/PmdKZ6ugGwQMjjxL1jwclCPSGyRBj9KyqkSbmJ5SShV4UW2
n7tEpwvlbM20G8KewgWE4OIug42jcJpp8nLnylMvOfPZqBs9e29NP4PEivwaNcli
xf5i0lXi5MM+NQ7oG0QAW8T4r2xzZ4Icdge/TAT4ffJPBd1zEDvRVAIXGmQvdSK/
iOeokIkKAa6KwejkIjUcFWTN3X02zc/jvJ/NhZUoUcA5YMl+sJOA8PPvVUnPSkCa
w0O7UhsFCUCB9OXQCsDUKpZG/6AZHFoAQMbK+gFedSpx3F/HeOQX4heAezlzh+NT
oLc+1LaNoWahHCBDC94kHWNOM1NBS0z4q8SDIGdI8MlZtwkUYHrrC9PEQ9M+aGSD
QTDntogxjHx2mqzam35VBdUe5Gc0ioztcWYmeyWSpVM6TrAlriWT/GihJH/1GqGp
COXpPW4ho/2TI1+EWiQEY/o/JHN32uDbUDL6K8e1TNzjzDPTTKL5yW0tKpC1xmea
Es7p9Wy1mFNrUwpn5/EnNrB3vL/n0YXjn+RrfBcO8IzULKaCbGtBsqyhQk+OimM9
QTlkfDloahbEEhdi2q+3A4jQLh6Q/+NZ+FQ1vFQ1+bsnvlkBO3EH68mPjANJKSFB
H6bGmOfDGzwxZ1n3WElLwHrJzuEvLPYRAG2beVvI+8EbRGxNvLICrwDnGB6aRbGv
ah0/B36dbHo6cpoXZyK55c53GuWHeq/cxV2AS8IQCo2zQ7dKc9o119LRVWAJhNFm
Vek/Pq370dPvZsbWpM4sOPs6RIqLOJ9bII3obr8ICxtbUaLKEhLyvOQGsquAiXN1
WKB4PSl32Ch7kuOsSvq12KR3hLzmWF79VQVFxqEqcxZIoGmzODM9fWGveX7O75Lj
6bNgaZ22BCtSrZ4WWN0MqUV369M0igMIe1XF+L5neZbXkWijB+phH+ooHfZduZ0Y
j40Bqzs5N5YvvM8yfjZOiuKojt0Iuguks0Z/qP7y/zwqAYtCMWPeHlFTxBrP0E97
uR6eyXda+5x3bmRPevwKTYL0j2+YOkaiP+OI5EscLGfB63h4CyodUQF58lrSC1yN
STs1ii1ie7jOQsktgT75H3eA6Mrqhs7xrTMiwY2tc9oLpiUClOH8SZ6tMJYYVs8E
qMryULBlUFFzr1/prrCIGnCs3zYGN0WcrlaUYn8L/mKyYUT7GmmegnJNzuDGDxlL
hN7oxCirUl+2d8er+FLw96UiRjpWj5H2QFGQAZxq/BoLw4AkDuj4XRbLCDK5PK9q
DDzmTXmwxjWlGRovBAk+2XRvc/FV1wHXOy1sIvW7GXD4qsVTAUAPGbn5ukfhF2Bt
DXBE/JdAz1+J6g4s+4TC2rhHKtMMBpLfu2h6ZZuc9ycbqeZHNsZQJGHZ6MBasHtD
QmMIBmJrXnooXw/qMEm1vtwyhCNECcDLWWcPdZSB2X2acBfGz/yxL+A/MjP5/Av8
lmlySQXNbP+A+qthd5gZgv6JY6JDOZHB4IM5YcSY0Bjm2+w4vMBbQa5gVPCjPphc
ejuie5YL04vNNNR5/ZKpRgEL6ngMNdFwYyIrccex5qbJfbxnIgKfbtSDY2giU/k2
ir3B1ne8vgScPJyLhZqw2AOQqGgtU+XXcquB9L2lsy+LQdMexoPlGvZwrpnYeOJq
2PEPey9pYnr5Sg8eUOWgM5qFBa5UIvE6XfkdwmRxqExNZv226O/qvhDRvm8r8ITe
i7exLZVN4xWY9HBU1oS0w/wsp3ZhvfcCmfhHvvOZl5qD1WKM8ElFNN9fP0oY1hxj
qWXYPruwgUXB3p4JCGZrETKgyDASJBU1iQDxV8OmsAk9gzt12wPcwA/XrwwPtB+O
ktLeCgmBl8wCWCd8RFOSlNd+FcI+NxpcPtQkuPJJA/egaYHuVlWmwci7yupbau0x
NaP42iV6MAA9ZeDElueKK2NZXQD8ebAPF+o9N1H/uCWg9X/zPIEV+ocb0H5crCq+
Z35PzV6WdSbLtpEWY7zGa5tTl8T5yUT1FCNhySlvs1j8CmQM074OAaSm/bEsxbVo
tTo2ujll2wG0pFrx0h0HS0Vl+0dG4k1qkz6XDN/X85qCuTx1lRZ0G582oXkXTH2w
7YZH7OEhyZe08HGEnrvDHu2lJQPSx4WM1/vnluMfb3ffjlzH4IgHlWQSi96U/0nL
wUONIzliv1d41tDm532h/DTsmdArg/gIcgPGptX57IMlR/4TAhbCF/sq4GFuBba2
eZRfgVEYllRXJ9yZHP4W9+yigqCBkfIGDVQe/Q8jTSkXeHnG2WqY0fKpfClmGs84
9ezfCXBI7bFhEghqpsOLfAb1Jx3A0TkgJ8sVpfeZZzqtNmKoxG/0nzA8Ay0AUg3b
Hd6NvN/W7GyO7QXov/aNc+heWxgA1fT7d7fEjXBjZAM8v+xTMymDWhf1t1eJxS0n
ErwTNGXs3uKAw0rFvIdYAJNGKhVl9/aziEP/zAOf2OwrVzOed17zNQ2UVd8p2YSm
z30r14z7HVcckYuwMV/Cx+fgNtFMgerS3TS8nrmjOL4/hgaIpdyuhlgRzmYI8lr2
owCvGgLpa/+jAkYc3CVH2e6MhK7stndtEDH63qjlMWRXTn5YWmFRrckOXuJeIEfo
g2Z/kZ5/SEQX/peFY3rsudRW8YHkJ29Vx609zOvxXKfV/VLQZRWhO+KOYWgktbv+
i1iptEBkE/Fhf1s2Hutz1Q==
`pragma protect end_protected

`endif // `ifndef _VSL_SBLITE_SV_


