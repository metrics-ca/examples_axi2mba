//----------------------------------------------------------------------
/**
 * @file vf_scn_data.sv
 * @brief Defines VF scenario data class.
 */
/*
 * Copyright (C) 2010-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_SCN_DATA_SV_
`define _VF_SCN_DATA_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
ZqHAl9MFyqvhUqnaw3Mk1/67YIQuGPH86dP3A7wOuJFZ/vT53hR0penNw4ffl9ex
PyTh6EmgcLG7WeAXhDz6UK3uEukuMf9zi7DUGo0694tGXxW/m5Rnk5xre47oNLDY
DoaIFw3Hnti9AX2RH82bTW1tdkvPzdHnWQFIMi2Tkgrpp+uXAH1WGHqI+btZ0U72
f17W98yqYSIwNYGjkBbnYAOylDtY9aw9RJIEHah6WbcpMOjK3Nv/nBzH5nt2KtCz
H6PNWzZeJxshiq8MIu22/1xTFjGJRuwW8D886dMoceftvyiZUqlkP78kLnyxKRDh
Wui941yYCsnc1ps5w91cjw==
`pragma protect data_block
T0uccK5OCH49s/Nem8KNF64f5qMFVdJfbTg4JpfgU1kEKh5ipF1ni4/3YOlbm2aL
zCckKedn6ddwEM9cx2Eue+YqDO9Sm1legO0tdzMK0NQSYvJ9eMiDP7hfNfVv8Id4
3akUzJUBbaP/Avft1VDPjiotn6Wp+eF5Z/ATugDi3Ag3DKa3X6arLZusdpaWoJ09
wq8fF7zpmoFrQ7taUo5fcLYczmAjUTM6Qz8jf8l5z+gWvyEMS3P+fukHMy4jkUfn
MiQm6RRzvGo+R+y6jj5xm0lnIdPosvARynsvT9Gnwhc4uc9FRsb6+vkQ7Fo3eKB5
hMTq+ednB+cVo9RfzhY4UyEmfkfhT8gFZ44YqSC9PYoxXnNMq5zXG0253JwW+OvW
PBU5K69N489jOI7MjgvrsU1opI785mTOXBZANOf0jSw/eeDm4KPghIgyATdphGca
qmDqBVptGVPVMciFxXPbaKfyR8SiNCqpqrq08fZNcjbbAy8H4h1VY17ZDZvuVmaw
TPA4fGgzYYQoNXxmk9fKHW8CDafZlkl/mWsjiJhXQCyMH3uBZ5izQ2WEuUf0g+a7
DC7HGFt+YhbivuTLLvwgI/SJkhXRdPw2+3FQCUwKxPKMUd6QuLKOREY2NlI1hYMX
BcLXPG9LEebCZRu9qZn9qbAs4x69wk01vz44Qhx1daCahdqEsa30IKecOovLJVOQ
RHDTQO620UXBZFMQr9w16dcvXd519lZGksiNnqpM1fiW0ujlTRlrZYtMHlquXJaz
Mj3hM5V2gKA03/EKpPf/wNqrhCCjX28a04mGgtNLfKr44d5eH+uxQrlQOuY8Mc54
YIumRZUegfU8dpMFoh5ghEtN6g2ibH8H1DPhHZ5EQrrtN9JQtc4GV26Goh9J0pXS
yORx3a4sE8zkzVHswsxhFvWXZSeE4f0O6J5naXoDfp7n5I6lN4ouHD/KlvX/UXIN
gwOg//PcTaUQSOYavSRVlCreEJU44wHe0RuiHJX/RjrE9JBo3/dpvHqfGxuldcYy
eOu4hLk00zIDORacRRPxl6j/lLZynobBldbzbj0huIwi6ObZ0aBGBoZfWWOjB1Mt
BgQ8crkZU4k6NF7hzxeN9PrdlWiomzt25t8he23Pa4YYSYwikOWl8hptglGd+1ld
J7EYmzdu4m9eKGnpk9yikhXlOhuu0s9WwHWmdykYcoICuA2Tn4SGbL0E3E2sWpNE
09CAAcfo/Tmc4RLbcklrhew72rUXIcr5wW4WkT5mWO3cddI55uSyPZODT2SSJvWA
nOXF/H18rUXsHk0GwodHwCvx6a7C3l+Ddveh2713eYHCUwto3/SHe0JkgXNqq8Cy
iz0oJV5H1PIbN5MKryouKgXoL+dbPFvcD+aV4mVCdktoRe5nJUHenuEBV7kQSEx1
CPyagZ9cGpMwpVmi6v1NKMY2ohGdwyHlfLCwFmvrspaKSkomcWsmOOBniI3stNJF
I/ByaMXgkvwzJfKPS1U0xg7WFBQzAcFNMd4AVWyPzOBKIl7Fm7O4+BnyH9mggxKN
Fqz3vqY547b/ixSfNAkZ5D2E2BMeNoXwmIz7jOWIiHm2s7k8r7p23QljyWZ9M+fo
iB3axGVFpDjykErlqbMjv4EhwWg1o3ZOAIGPcpLoMvkzU5TKPt2nvX7XBNSG1H2V
tY3RMhC14N9WIf1W1kUOjoPROy0526e31ILfCnu2NC9a3LHewH0GmbGYHmznZ2i1
+3TJB/4294lBMYzr6P9Hxn0h3WuQtylJOwPNfUwHBzlfXnKl3S1ByFa/5pvQC/Wq
99RqOzItYJEWGPvYyfYaUgHnSucVGvKqC/UTyVl9/77xvC0Sg7bRJp+wlcfvGZxm
gUP9X3BppgdfFIPFFPjDYexGhlTDXKyEs76ZpnTzGn53SZ7QvTMSdGCp+yrHLn8O
tkAc1LMg7yy4y0PT1L3O0zahKUPL71QeE09xTcPizLE7mZL6fqcfrM65U8bF9DTV
c8b1pue2alLQm3re/STT3eUHObbHq/47TLTTEcSRfbnVO2kUuhacSsVSWPycEFm0
tICNaiKDjkdcF6n9lUj80MFEdAo8G2KLXOAZz0o8k95Yp+a2J1G5qAsBizcGRFhN
cwFVtekjJUzKTbHQdYb6j/aUZbs90oq8IABNlkgPNE29/U+nZ5c0qok2/nJpd/yZ
WXkQH/RmnxXos19vUTCaB3P8LdUuBXJwgbaNf6YThCqRQXOAYeGDlYvTgTHSQ5U2
unTuoxEgfybMNlgj3LSmr3SiomWvbudXoM/Z8qfLR6JrovMFlHneb0OLNsmvQjIM
RZGqKcQgwZBh8VvkZ36PJ0AmcstB4kFsmP+IKDXbBDXg+fy5lVxpUkxjYlYwV/t/
arsAVCtB2Mmi0ZsYQ0F8ZsS/yizA9SjDMZCiFRvpv7Is112GeFlVBMXBHeMFO8iC
Cl8Kl2bb2zkpl0rsUdAt/XXBAYUE5vEJS6EGtK0+IrPWZUxNcWrj4ye0X0b+zoKT
4VwXU8gPEN5whvwKs1ydmPcUwMoH1TBtfkgHsa2ZETnPhV6PfY4/xp3X27jvdvJ1
7qMmJcT47AWNcGnW4ug9LMOq7KZv4TOA9T8bSvexSEyECJPyFnrrJYNLpAQ1BAHs
nuH5K3E6vRRYw7KOuaRgbwReK/CM9Y6MIY7+mq1Xqu85+Ls/J0O1tVFvN75Y6DBH
/oQXp/WY22dhkJB5sMMZ91Mha+vMMsww5m5g2Z9zPOt+xBrSnoJgMIjhbfhKKucD
4zB4xzKy96ciK6iWt4CPaXIg18tfohNPYbgC2UR6BfoXG6lQjZgl4srNyZ2tBqGs
BNAeZ6GptDSg9nPLdp0+FjIOFrE9tBnpyn+mGOG75MTEGj+Cn4z5PNPbvJ6px/+9
Ni1yIPwX0Duwe55Fw9daM3XITKH4XEDR/ozPBK98voxK9QYylUaRC3jDZbWlIGYG
ClI/5YpmB2q9d1n5jPfl6mmkL+kYVmY1PdOjrYvaBBwyr7HKvPAI4hDEd19pE1Ma
uo2f5E4fdjPY+FhUgS3Fr/a6IabfmzKEGaJEZt2BgZ2sNV3Dgq2JEuuAhn4yqeHI
a8JBzqIGJIgGTacoZIje/sSkM6QqWGWMYD1B/fgmOvQkLdPFyWh8V0gcapPGY8ET
ozLAU9IrpVUqxZHtt6hhZe40APdzRB/V2hg/CquUTmoDNBLB862O9UZVbLg93X3v
/42OT9sylwu6VYdAfuVdaeKnxogVps/350+JTEC4VWqOMoCzDJPSSNoOFSj1hmUB
79ADQ3xldCwkGkVDu9SuGmxOIuIYnhyWH5AnVxb9+e+TuNOJh8gD6NmDIVeafcri
RP04EFGrvOytZsYWYB3rpEWO7e1b838cZhI9BTxeclEokD5EvfqKxb07PEtHR6t7
iLSTHUwnk3Vt5meIU3lsSlhf7e6NTu2wKd+S3fBIHbcY6jvXql6gnst7EmInoExZ
6zxKIO1QFqJo78yBpQvBqZ4LuwH8Rr2qGnPHDe4c3HmexDitN1x2y9Rf0q2FblLd
awamvgSKf1s/RzrvseLrfPno88+uSshhPCSGGv/VIl/pyYrRf8l5wdxb26q0GTWe
IseEpQQBg0aIlx3za6KRkDLM1+Ni+3+Nv+b8KjdBiIDb35ZYyxqqOuiDushaEbfi
/kNRh1cDloBrHvU57k1B4GzbpvU5e8YUwSBGD3Dylx/bcUeROXyOAnUv7N1dhbJ+
B3XZ/TdjopU9a0yIIyLuzLbJjJgDqNLdYoFfwv+0Hi7EhyHnopACo8YkFcFArIhF
BFgjWkv0f9NtN9sycbZXv+5UVcgOix9p/oWPiMpRdyBUGl1daTzSVs11vwvr3OYu
tU1Nf29tdCqr1q9SZlYSm++j70DmlnVr0pXuRhic/87PotNBuUczBMBNXYwm2aHd
KMCTB04A3vV6SHZW9tzBVLv576HryFpjJoRgba60hDniSIJwF0+Xn1+BbX0e4CNB
pDOcv/g+YTomsatxHPRYCMN2g+HPhtrTQa+lv5GZZwy9BinRek8+XhSkf7Upn4c3
e7UpgLprx24C5VXaA6pjDSaEB0j+jff93+HfbwWJE+qV3B724m34ab/suB35ugWt
iWjjfZOn9LPyq1SMOGV7jbceXA8B0FC3Ps8v7GfLQnfaq8nD4AJnfR1eZR/hDFNS
+iXYP4JepakNEgQhMuqyXXWKKXhrtwyf4tpxShUlB6O8d4mTGo8EWNPtTzy3oYT6
kIaMB0KTUU/J7AIImXqm513vyknV1rMoO8+huLpK21PDaiKIWX5RANhJXiaZvwEc
6eH3I/LDUUpLju5Vs9A9nZZmWpfO9nCl1mxjueM/HXRgfnMByA3FaJJ88zXW50Ur
L3rT8eLW2X2vR4HXbt8qv/v/IsTo9r1xhtEgGghSHwzc4FTAN9fsVrCdizRtH9RY
WFEVAYtvWqggzRHJKZs56FJk3ZsSAizK9zPdBo+CdcA9IuoC/3l9joWVZa7qpS4T
p9GAJwNyuo4YLElxPKuVLruA8am+ZGtuu+D/K6KY3Gxk15tIcOSgUXrcnO+QQyCq
WoJ+Ymqw7S6QJwQ8/4y6xwV1cVe0D3TUAOdPD+ymcH2DcOKvORTl5lioZxkBC+SS
uVF7Wnf4xNgcebgWJAcm+hRyDhTrIt1oJlrxrzTbnDKKfonWVL8XRpvEfOTbDudd
uwC7CpFw3cOPtccIBrWWs4FSEuPrdHxE5qE7qKkVPaVsNWlb0vPNd3AvSbXj44f3
dGH9aAUcnXMG5GASj60Cz6oBkm/+QNZf1mhfUrh1L9Gp8D0gN6bgZMZaO7zCoi+W
DIcTNnG6OU1HhBHj4jdHNXEsVvFXgDkJq2arRO17GM8j35K54g441eItcmC/M589
iGjbaF7p/nWQh3M3aJLdLIjT7w1kavlVtCiKMSIBICrjqnKInSHD3Oyy/odraA5T
9cVHdWcTyhb0fbBkwrZSmodx/FP9PQbXTQaC9bjoCmdL7VuuvfOdv5mkxgjuirSw
FN/+XhOhHdi59eErqnPZKnNpAnkp6lWpnjDz9nlAdeF4i0rk0FSWCiYz1Ru34e+Z
idRj3IqvB4u7YtrNt4gbw0dK0rm98udFR6R+hbLSeVUVXjuJqZUYkq+CERHgkgdJ
ZIuKkHm0aKVFi0t/B+sP4hj8IVDKjgnPL7YSnWNmAbArWH0pOaymlwzMJuQlPYrv
jjWsiNLjTNU9lqwGBA/rKnp7STfVSPIStaRdO5C1EHETjS+ZwsuHmAK73iPJPhZN
5HyC2RhB1vXFqQUP/L0JFNa36/vRrVqdAqNrXaJN3rtTP5ZNoa2dzdfUTJm2cxEm
ShD+jpAUUDPgKmvbSz44pzEPD5ESy8PWwrh3TMQN4Z3xTYs3WFEpA8cWOXkH83/k
V+WJP8wse7DTqKeWXF6gFnUEwo0mi0vnV4vFnxydMZmStDvA23ykl53Ry9S3mcjz
w5FRnNkDr2vh/JVfoSL/O5N89oQeyuB+H6lKG8CnCXEPPzXVEspC7iAJvy9Ffvbs
Q0dnnhWHft06JUmpSzC/hSC/3i3CeIPh+7imnzsdSQWFUWiSvvzatYnvaMThQVT1
S374QsbSbWf+dsVYu8HyJW8G5AqLDmZdej+2zOAFxMi5maxlocSHwAAOI5p+Xmut
KsFWGh/xNdfFksfyo4psPqFZ8ywI4lblAfcc7sGYLpfp1vkREPZ/a/R0/IN78mHX
z66ZL74Acbgl1TCMOP7ufJoVRo16b+3kaTGIv9RYKtGCVpz6x/qG3zCOxd8OyEkx
R+imcAcizkRbxjeskslQ4+BabOTU6i8fQaQ9uhx2z9i/aGyQgIW7MxI4PHsh7PoW
kHZvEOUR/8modnhufOJFuBHGXaKNK8Hua/M5px5PkIWkR7kwUTvl+cdI2wbUJ7nI
pLGxwaLh+tJ3yWWpXal7BMZhHJ2RvkCXkGc8fiFHXfw0SQlzwVRAydNt7gzJKRyA
kqC2TkS9dktJN3JzFeL045Cxh3O0HG7vwXvR9a6NmkCxvrz91qyDhAO4ahymdIEW
uUUYBeQc/C28bvfwdt8i2ASWX30c/TkWbP+knFkmRQlJoZNIJ0FjlmQLIAkOnPPp
UddnYretCE/2NnXUYuFn7hTOT1MaizLTMJuMUEVxhgGiuuX9Uz3RAkDby5lUlwGV
16kcl0dEKYPRXvXuQtXXmG4NHATZAAZ+qnKiripZmLBTOgMrKRbqwbsWFmbRoYjs
Phv0ByDEXEdqZc92NEiuN704tgLqzRo6u/JbZvYPsLJ4+puZ/1gfeWq993bebMAE
respy1AQub3kO3yJf++1VbBzwzICCvnb9eKRxKH1FtY9MbATutEyts2sktpvWKTO
9cJY29w5f83LkZLKsb5yxJTVli5Rf8/YVp0MM4q9hVi7HzrMGxn6tQLys7PFGhKO
DDbvo5/1n9PsyzwGwEesiW+88r9rCLfUg1Mic2LfnrTEC0r1L+4cGEq2m8U6NBHm
TduhsFOH5Qf8Z02b0m3ltVMqRzwrCNXq6NOJHZBhCX7f4dmAPT6b54U05fpqN7NE
gYgmk1+QjdRIleStxjNgX9hFdO7aPkgjgrZb37Zlno8AJJI9m3mArXcJXmdSfJoX
FlskaDHCyq3JtuFnpku2JwHB3u0VfAq++98HQu2RENTxkID0KepAOqEO606W+Obq
wrbFCOA4JRDm9TTqNxjjHLBXVM7Q5y+Q0QNTcd+JmkFSYtay4PJ7ppF23TRCKY7G
DTbGzYAKyrcwtbRlf0P9jT1NJMaFuDBqB2ZKPUIl821vvGBXXIYkNAoklc9fsOOG
MUPLVjnUsSta9zJ34dL4bwdkZOMbU1DuZ7S1tsxY1nNIBHaZM1TNLKWy5KhfDvGb
Nv/MW8lYL62u8W5WNURfKouyZd0c5AkOHmoXc2+UbqKtcJg9FafS79pvfRe0R9Fd
8YRdVstdkpAT/+esO8X6mpv4sV+29+PZKH4GXu4grni8ObG+mXmeBdWOHCPP3oRu
9gCAMca3M1WGkAp/Ksg5ZjKhNnvzupvPoye0Ud7bjHeYTgG3zrOCgIeyuiHwsYPc
rFw7YL9b+lmMfGUKDa25n0sUVAaDD6sGHxxrXjgq/wSPB4DvfUztyUjnYoZ4LktB
sJsC8YfxIDjysE3DQyF6pY5IK0L4AzjX0duEJCWrqcPvZxmdnwlXJvuIyAI8sYh3
2NVgaVUxWskhCDrw0iw5ZY1m2tR1LJXv+X/EkLP8C6U3/w8uHwGGTYoWhhd7TKvT
6echF4/szCxg29F6JQVe4urNMOgaBzfarlXLa/WNWSUPMj3aYhFROUD/eO873YmX
VLynW9akD05EDMd301mNqB2/TtG88u041nCU5iMWfhE7oTIciyl9QHxdnzFOu/Rq
F4NY6lP9nQ1gBzFXuykmy0nT5UlIT7u89RdnOKNRV0NVH9EAlWD4eR1ixuQGovZU
c9HiTuLtvY2Tv5migPq3Fhg5zXDJtcl/2f81JV5sB5x+THR1Lr4bSdXCgPLaWHnF
MegGOheQ1lhu9cUx/ZmVLHqnqE7MWuZh4p+PXZdWy9+1hNCZD01tyPj5XuLGZl+a
a3sayald3EtMvh2HqXsS8gi0UmiH0I/+NHN7rUA3S9fWIhtJ68jnunOs/c4ndc0Q
D3hodmilKjI7NeZaoXkQPsl4KH2t3qkU+l3qfqyeb9kwe9DhfAgzLYCn8Euyxaj+
QYcv1C2gUE//KxR6SWiRlAJcs8PE/4/SQQPMSVrawbcSDqeflsNINwzk1S8Ozmbz
qkwCZjZvaI99UpPd3iPxZJj1lb3SoT4iGs9hM2QBVTiOKnsP6b3fjOHaJ5W1F9dr
GXOdPpmzMqRhGhcjUGtSIX/dBAh/8oRn4yKbf5RVt66jjGEmTX4Zlrv96sjc9D5y
pO9xZBYGQOYBEzUE8fVr1p0k1GVN19CkE8jHaj3s9bPxofDOKFp754kGKEugXA7c
dXnilMhR5snEyH7t6e0HaffdPDs8s/dJ/ObmbuY5Vw3RAtvnO9WOQu2tfcAiCK08
qSxxavKl2fqgA+aNa3RX1R0QpZ59pB8ACRf10mtkmcZYSGlLtsZZg0vVuNqPD/CA
4kT9U/XdwqbzlTXho8VmlzuJk4jgsSDZGjF91owhI04is0+R6n8WZSl6j5h28RPr
dBTx/XUkFHa0Uo07em++Rm0U/QJfZGoLZ/l41DbIMgLS0wEIW1mBOpS6Yv+e4C/4
vKYenC8NdzIBt84l2dKGugzqAK5urtmf0NQ75oD/qEt/lCAzF6DvD2c6hHeqKnEd
TYrPNcu6Vwoqf3G847T6SjVdaUQbLIw3jg7SXnZoWaVVRjBmN2wxYH/Q94TwkaDa
7lNYpdBAq7yaBzBuJ6Qy1YXiBtp+8aRSa13Z5gldr1I9yREkw4aWg6hXM9hKqTUf
wpXMRrm4AAYBnw1ifKCyUCKhGLOz1Jx0c9k9BYq/PXlTOpSaWKYLWGCw8BBoNC9M
rlrs0wAWwRJFSP4G3JQL7HVb/YX6HufeyHFYYvuXuQyNNMEcq3dTpTRWmvC5BnHJ
HnhS5oWi2XXSY+e/Rgod+2uU7nvjZiiScGaN6nyjtCe6jpvJL8SCLIRAkqytcBS+
l/wiCoGVVqmXXkGKAn8YWUXesDaFLdyu+3uzhfY1bgrYTuyx5+BSUgN04tjroXQq
IhUFt0pVJTpTrJ7P7eld7ij2RNGq1sIp69TstjrTclh6TRkJUtinvAC7/kHscsYR
Rn/Tys+kzeNzb63/LsKYdFhfNsnwbqCpU7gPYWgInjP6gIzS1mEEGkPtwfMTUlE0
Lax2jjezbFgU+9cnBhN4mfdNxuMwgGwaM0wTdBK1K1vCszSctkgOd+pA8AjpkM5v
r7QQAO6578B6orFR+jDt6sF2uLJtaGRFaWlDF0lYN3pF1LHJAC2U1T/uxun6rU0L
fMa0FOrKIG8ZOcB1hndi4gdXen7TQmFfPlDqWl0I3qCgpk70zXJeyd/iO7AGZl2C
NRtbEZOd/dmIilrDFvux5PdL6r6LX7CKJ4XVI3MbwKC4LOLMtFiNn6Hp+8djgs+w
Ibq2z0pcRNnX5bVM6kyvb8YcahcrvwzRf9TCbZI3Lcejb8+RhU0K5N6pXsUMlzel
E9Jvi7q9HafkpHflW/tCLQgRXNNuC23uoQfvH72clw+Eg0ZlGD8l2kNTpOpqaDxG
Y1W3FTjrOgBYHlLB9cILX/5AVmpV7OVIF4fZT7vOFL0AzCjezlIGUpn6APXnjTGW
0MKzPT+n99Rkd2vIyPm5OIh5kOVuHNVutyhJwnOZcQw0VMQGNu5nUG817u3fD7In
9sQDRvN0Tz5IX6137MU9bp1wiYE10AtfeLE98gyUSYIgmtlaTP2h25vve00/NXxF
jCRDn72WdaqlGdYfmCzFGlhDUFC6DOsJZJ2WPjJi24md233LCzFoTQktudflu6oC
JIWyI6JeuJYVEZPUspjB+3eSaBDnN1OtSHkaOZacId4eWYcoUtbetYKewJBLON3v
Fc2U1kWdnmeSlbrTQo1jELVRwAAjrya7CZuaiUvTLUJ1UCArE2bxVo7tcd2XmPE6
U44n6B6dhUSYupg5lcJJvknlYPqwMgmzNLo3KMfA56R5tUyZOxduqpP7s6C2Qjuq
YTpo7AmDqRVzncZZ+9WNEqJkixODWO9vJO+GShtRJstuHfUAdh45fzJpt2FVE3J+
WdL5fyFgMlSoa/Z1/7/T2ashQUFMXcolQPRskq1EOGcox2dH74CdUsJr0a9Q/k7B
7Tz+wIHxYVjS5gGI5kTvHmW+T+J6XGV2lLBTrvg0B86qoF/xvEOfAfY1aUzJfS+V
MQ9o+/9saHLRVEKW5FLY44gjJgIkVooN6BeEV0RJ7NAId+3k1xoE67mAdiuw/z4P
lYEw/LGVlV/VBmoHdfkYiSZfrnM0trenlTzgCyg6OSTs71Xi/tRjf+FpYECLKrT6
8CTMuxNDnPtWu5Ou5I1TaaAqdQSh5PTFKE9eYj9Udh72X1cA6r5KOVYQdCv043mA
rhpFkhalGE4Tffl6A3wQdeGwUdHFUCuvsdn02yowti6CaIvGQDOPfJW20N+MsGrn
k3z5gvEaD0WbD1DFCy7lGbyMymIgacyzJycz1nNJjlkASVEJX8vjMYd8I7geLCR2
qc11Ezeeccn8XWuewLSF5fnrdwg0wUQFqWyxx+Sh7A0px0SaKFEdx50JgmOKrMxz
v1/4pbIBCAD5mcXX429m42Wg0UdpfWvDOg9UpjDGDO5bSLDdZ4dbXRSB83VgTpoV
OZUqFB3CQJmy4cMyelhTY4+eg9KkMw5v7nKa+vpqGfWy7Vafh3vYLQZzZ6/A3nfs
lnrNMAYw+Rxw5fatDITJVQgHTcxIgUEAi6CCgx7wc0WgePPydBH8VKzIHT2CqSz/
3y2LYBIex+cTUFjMP+UrliGp9TSHcb41wIoHFBXZhF2QocCEPUzUxyPo10de+mey
nGbCYTzzLICNQ+4aDAJ8Ttuh6cIKeFngu/Sy5rQYivFBzdTcJY+m0V3XEYIxQIek
ZTh/9KbIe3/J1gS0wBOE4zhQaGEgdjuracHVnLNnCL6SsC5eYX3JNlgWtMRFzF9R
c9qQaFdGtn8HqaeBhbS/EePjci5RfRXIIHCyrF+vJFlRG+7TH6pOxWaTWAecBhsl
5/6RHo/Jx7i7mx9CbwJMm/QA43OZNTsTtGqH24wDfqrvS4D8S1vsaNa8cMDjNrTN
OVUfRGNykbNO7TmeqDtMHDlBtUqr//jHxg1/SUSrYt4tWeEP9b/jo2scR74Fg7pu
BXVOP4woMPj4iLAcMW35o9Wl1NOk01S6bs2fQrgRWqIKzOf6XtZEEzVmrsAKn7+b
XX2kpL65CE6EFN0s15e7W2174EzG4v1qHymGo6aIB2ZLpyDJvj3blU1g2Ks1OQR7
G0Z/h65gwDGkHFvEkdUlY4bh16l1WRjboGdsTBXX2gzlFnJI3Zu5Pi64OqaXrAST
ZlhmHtMpTpTEoWp7gkBU1nKj6mapeuEEUuUpOMHSz3SvUFA7qg0xpbuwY/kn+IeI
SgjOOuReHIuysi3tz1NjkA4mBk+3dCUCJ2MntylwkuUelslTdKiakE2G81T81LBD
6I7EBXTc7QOPQI8BAJvvNS5yfasesxbiVUYkXe0T0z7d5AhcGsFWq3st1iP//qrT
/bmi057YdYVS+ds0m3A2FzMaUQZk1+Us71OgQpf/DlTpr6/QIym3ljTlUDz0m3rd
rVagNVaklGm+qxWMHmHqM9m1JZyPiX+2tAcLJPlKCNo=
`pragma protect end_protected

`endif // `ifndef _VF_SCN_DATA_SV_


