//----------------------------------------------------------------------
/**
 * @file DDR_A2M_ADDRMASK.v
 * @brief Defines AXI to MBA bridge: Address mask module.
 */
//----------------------------------------------------------------------

module DDR_A2M_ADDRMASK
   (
      AXSIZE      ,   // i
      MASK        //, // o
   );

   //===================================================================
   // parameters
   //===================================================================

   `include       "DDR_A2M_AXI_PARAM.vh"

   //===================================================================
   // ports
   //===================================================================

   input    [  2:0]        AXSIZE      ;
   output   [  7:0]        MASK        ;

   //===================================================================
   // signals
   //===================================================================

   reg      [  7:0]        addr_en     ; // combinational

   //===================================================================
   // logic
   //===================================================================

   assign   MASK  =  addr_en;

   always @*
      case ( AXSIZE )
         P_ASIZE_2   :  addr_en  <= { {7{1'b1}}, {1{1'b0}} };
         P_ASIZE_4   :  addr_en  <= { {6{1'b1}}, {2{1'b0}} };
         P_ASIZE_8   :  addr_en  <= { {5{1'b1}}, {3{1'b0}} };
         P_ASIZE_16  :  addr_en  <= { {4{1'b1}}, {4{1'b0}} };
         default     :  addr_en  <=   {8{1'b1}};
      endcase // case ( AXSIZE )

endmodule
// end of file
