//----------------------------------------------------------------------
/**
 * @file vf_axi_slv.sv
 * @brief Defines VF AXI slave class.
 */
/*
 * Copyright (C) 2007-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_AXI_SLV_SV_
`define _VF_AXI_SLV_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
V+6a/adu0lG9GZ/9VRomjbvL4+mNxR2h41dGocwS6+Q+d25Cc/7XkqNRWjgm7psp
FBUQ+l2+yecuhFmbQbXhMbl7QkLCB4P0cEA4LoWdr3Y/VPlEG3Df5G81snZn/Czu
TosXbqfPlZ1iRt/FNuHpWQxoE/OYtdQkVmu9+twECtTplLZlbDO/9Wegu/n81WBo
voyEbtks5XJaxkesltUTpUzflRWhR+u+zOlqxIKBoCsGOQKLAVHcTMsrPL1UyZ3H
lhw/qCtb64LtI2Mzc8qCf8aS6R1XFBfZ71IcJJHmpbcoT21pq9VQlEI1dHL/NGoW
PbBZG5CuJwYurry9MyvVNg==
`pragma protect data_block
qzOhL4HW2kMxY8ecrdUQjwkVmgbSqhlUVCeGzMI1c96KGUptKAFwm4/onjtMh14i
NqvsdbqG1gQV+SBLhn71HQ/RYkK3G4QDwt2C0GqUwNdcCzcHYzKMsZ95Sut3T1el
d60DsWFkrBIDbJR7h3QqhTbCIfcqZ5PkDhn2jrgbjp+xIXT7+7DUX1rkqdRT6gwd
X073FgXL4Js3bZ3wNl3vR3lVpkloDFjl6u+IeG5tzeV45Rlv8wIyhEtx/tfIEziv
w8ebZuJGmsviM3TjQ1zCPQbkNk7eioVLZc5dTwd4uVUz+f7Z798ijMtDwxRuXa0P
KKbxHl8bZ147l2TSePISGksWAvC4RyRfzrKmdHsS64QRg6CyiLiTa3ERCl+KtNno
jKRZARkivFTEcrqCfnekzWS/JayWJDI+3XLwuGDaIGm6vV5kYkNB3595PxALMk7O
Qx8wHJbbquu/6AW8QZbugrm1Sl+2Anuix5CfDYcL64HuNq58VlveZpRhFn8sFXYU
fokxpOXnTGOLIMcKw4UQYVsyQA1lINTW7UfAtMlDzdOd1kM6D6Fia02Z4GuRkIRF
YE/HOTe447/Iw3EAlCd3EN+fOYVU126x2G4xTfyen7VGLwxUaxYTAbDV4NNPOI31
uJA6FDICilfmA3RrRAdCNB+Or1ELOJC1F83bKtcldV24I9wL5e1rGYQk5bTAyLXJ
xqKDbEIbCRZYPy1xHwo5in3u7I5At8mUrVtLN61Xzk+H3y0/Y093RgsS16t0fvDN
I39znLZ0EnzIT921vvaHJs+aWaBazzZcIWeDiyjc79Wp7G3Q1/L+vd9YJRcbG6mH
N73/cFCQ3vxtC3wVCMqi71KQbXWd5Zg0gNgsir83VwN4h8NNKDoQod0e7q76AVW/
4uEGSrRw3Fe9JZw0yJ+2kzow4+2INfxcZB0nniXIbHoXcuDhxdL+IhTOvTJFKi/N
tL6GrBHG4HVO55AfuwhNJkGh4bc+X2frOQoh3Y+W+DlrgV9nxpOMqj8KdS7/R031
jyD89osBxbdkXSoO1GyWDFaKQ/F0Ys+7DOsXmC+uT7OlpqJAXAz6axJOirzL2PMI
uzxB6p07XCkvxGtdXeayOSv+DoS35Crzp3ptrKgwMvOvATwehD7ZPcPQEATXp1Rp
BJgHoCxFAgpjgShuQ0wgnr4j+0vIz1Sp7m2tkQuY+qCd57xI8W1NnfUJZKH5GDft
iQvsgptb9voMP4gNP/DNd3+//1WXlKqDHwI/ZpmDQli9SumkExbJDNKasrOfVRHj
bFBBzyYgJNxgaceBW/VAAWViIzaIbSLv2dre4AeD6shgnlOeSqvGCsDQQ6ljhGfC
KrTs3YYS2Qt/b2SaNn46xVaJ+pfZ5zTDIRH1FBATCRSfubjElk18JmWQO4nm7KUU
u2BPxAdsGcb7DBIZTzdQOf8nqjNwJZ/Kz7tiqniAhy3cEy2/3swMD0BgRqV7xpiJ
YkKpMS9RFM7UdBMAeLEaHcmbob5XajZ+nQj3nu7wZ8pNHPoLcmpaXbWdOSpULGGU
hmjDQ0OV2z6MmVnu3aK6c3k06BeW0xoFFnIEdDmrBfDtm1Fhqhb1Pd0yRQNkgdLn
KuV8EbKojREq0JLvCpkFM/Ua2iqpCZmfj8qJZaBmF4TBhDJywDDKqEh/ZczCz7tH
VdHNKPX7rsi7QBUROO3jfrqHoBDyNOtXuZHeiaotdxivv2txSWEx1tfHb1OWX2qZ
qLK28QutSMlcBhmmmIhsPqLvbpKWwVgclz1R6qIKYYDujnnH9lnl6P6LEQg8AiRo
IC5ivoaYoX/gPxjxxOqPBEPHJQzrFMzZhQEnWdvudDRgLlt8e4PFQLxc4aXvtfBC
63C2BQuGwF2LzOjHvDCiCOR0wlqEoV1uR4s+pcON3yKn6qMaC09Fmspj1DQGiaNW
G1OsF4UBbxKV5QSJzCg0zIL1JS09EmiigogrURwEfsqcJ1wVNn0rH1igygJveDOm
n885dVfs/Ty8iMeoOiGZSLt0mS7NHxErcQisL6tRBb+YrCYs86v8VDa6ZNIVxEAN
T5vljdKLDLEtNy4QgdYxJ6E8Zr3RpI6CSAlWeOx3ryqN/Ydf2WolqSdicC3EKDTS
4VhKERpH04zsjLu/GxT88wqJdMOChPpiwyCCT4Y+1nQaKpmUDBlR+sDvHOapluS3
zZORT7IhT9ucARtVFx5JLaXbAmYRLvy8xNcE8xPZO/yEkmCNHoyyP7TPYnj0Qig2
XeHsudu10Dpg2VeNxtDxatWcpQADH7NpBRCh/GdEBbeAOkjPVxqNO/Bd8ME7kji6
ZAflxaofsgbNMfRbm/klh/uwPsfOcE79URlYuuTT3QImBG/+h47KVbe+kIxjiFYi
/tBvundeb3dNEj8tJLwalfRrERFIwQR5UFCzS4Va7W/wNahbEeRTek1mUf81KOVl
c9OHiVmVB8cOycOITJXif3yvjDFTktOEsmxUicKSBcU0gx0JY/99YMJ9ijheDMVv
9LYbfyEpqVa+UuGrqCX18F72+rEV5dkFvaHRwy1wXgD7wIcPn1nDKhIhrtX1K2T2
R1g563yZIhgnvZorRAGNmA5IGaA22wyKftw0W2dba4UBq/YkrBBHtbY2etahO4/G
QDzdCLpBYIBOsTc1HLveAD4/C9t86b5QJQXlfJtCEvypHmyTq5lYmC7TaJXcZizP
ivzWmJ3+42ZQfBTLVPNjnMlj0Xh+c4JIE9FMtVP2asN8kAmg0yq8fJYZ1xYfiK70
l5KJTniSrTuozmzKVEk92DWi5dil9S1O88i8Wc8f8zNw3qIAzJ6MwYFbfcPV4l+E
zcoQCpAWHtdsw+qxEEAOOuKeC+xm0Wj5fhgRJUBJMxURgSNJP5ATBh5GK/aAndKe
lbYrk4DtSMAxG+BvY4fFWTTvl3eOLq4wJ41Od55+SvCjWTLEU2nWGs9IBc+qzjGF
UZ2225HbrwQCvfFxPr3S7qNGqNMByIsH9qqv3ydvKWqctYt5Taldlg27e4gcziwo
py6bT2FPyiGzh411Imwodesz9ewXnIZm5HpQI4mzRvvyh4MUVoVdAfamN2k/Zkt5
9WgdOtUqNuXdsYrIKUkQm7xaeKljI4uI6mtZ1jyls0tIcm7/+fMS7mTB3+Qeeff6
3KuIEqAkQ6O+VRd/BEszIROvnEtyqjnKeLcajY638M9+/MayVQdCdftk+BdVdja8
DJaYUlNX09p7HFcGec+0y9XBvea6vs0zkWRbKRvNIMCx8OfCCthfkxI3ONtHemhG
Nbm2BDIyg7UaoRavynRu7fVDUAeV/hewV4Qq1B4eLE7m3DuCPretwd47Xxpv9mgo
nnFBqShxRyCX7T6LbYvXLs/QNExLvHxGI5zyHD+KQj0X+tulUwAvWy2Auj4hjyqk
FQbITF44ykRiXf3JccQKcTi4yJeD8Gw64lC43a30ABRznEx3/mnFULz/TvUo3o8R
W3tJPRgxQjSByKsM+NhZC8Mq6zQJ5UuRpZ1EjY+a3YaoaPEE8tWy/p1ahPDsfujM
eVQQa7dulIKVXNQmCeIvIi+y4qQ1Diw2e2MH0XaOu6Teth9LJ19hF3nF+K2NAUI4
UwCAQnTOFG2efRA//xnhLhJHXNKg2m5M4MYrIb8lT0I2cnI/BfS7dJhuMe1NvB2+
yn9RAYUH86I0WjfHc5XLBom7AQXOhX5e5XuY5OjNa+WGH9GdLnaMZMW+9QVGuWve
qjdrYhhYLoxu/vwz1as9HUYG49iM3G8MBfrzhjjrO6uQEAIWzBwBnRK2AWyqKERb
eWuzsE22Tvx1KI++X/j7bUBlCPj2Tm03WSwrH7Y++VWbjvWRl5/R53ckb75v+oUX
rjURbOxQQFxtThxcT1CmMok0Rz4gO/3FvMitlNk70Dda1OM9L45wZagFnLDTbhOw
YR2m3/vnpkh/GnQS6U+w0reqJ+HqeB6Ai5PDrf9CWf7kCcmRn1UcdmGZfFj6oIwN
QJTfvniC3rCtbUkQ1347KUY6PxX3OX7OG+MXBSaBeP0rmUrEXP71B2x4S++1IRIM
3WevYwz34n2au88dqsYUf8WQvgYEA1ryuhFOPRTuEQtNjCyPTy4ZM83NsQ+sgLqn
OB2cSwS/QMRYxXcmBm65p4IfqLfRfKgh5VST9nS1pBGLncVI+wfnMwt/V4sO/9TE
sctHolSNEYK777H4f5em9c/t45zprEVpAFsyVuA55wDpnsV/URGccxsgwAGBlJwp
oqCh4M5AAyi9u5k3lwvxNhI3m+EET0t19v4NXLo/nHIQlzQuUl4VVtmpNfjTzCbz
mBA6+nnP3lSIy5fhcbKsIh3HG9EMCzyoStw1B48b1ssn/u6R25ycwLv5C5TQLtWK
OGxiNW98KiX+lk06S4sDXQ+kun4N4kM8iCtgyd9Lv65TzsswBT4Nyulj8Wf4DowL
0RAOd+G+IXStYcAc0Lif2y6e93w5YAhiljoBDdXiFWUKvoXlhhw1QPfZWLm5eke3
PxQt20zD8elB34h/ie7BJk0WU35tUTPbMhr+Kymb4nTSdb5+k0SQIDvJpbBKzCE3
KUYbDVfs3H61puZ/Fw6YouGKfYKU5Z7N1D78U8gZb2LLz3vavMdn2/ICCV8amOuI
jxCMe9z6eJMRhD1dyzTFz5TCt/A529fF6okhA2cqQUyI4bYYBgxrEKkK/k3x8eyQ
hsU85UtAUHj1N8tglPDdyjsq7xvE8325usEtbXULRYfx5Pv5cYtbJp6frh7nEBYj
div1nup94SvkklSq3AnaHIUJWNIpoxN2Pj4Bmo/TbDboVfo43tr1xB6Ajew0QnI0
GAyCWnwWzQqWxe1f06CDAM3B6tASmIstUifx0UBvl3fQc3Rs0w/VggCeDaneRm1N
y+fTbL84VrTp2IyUQjedNBEsA1Jq4uL5TMU5RMlnwgDc+Exoqwvm+T3GeVpj7eFN
4Pe7lzRTpTOCesSAzwHE7fxd7KjJa5VPbAA7fUFrw7QLkZ7/Ha7f2mh+MdHfajZp
jv2Y/3KaZUB2csTxx5FhskaylbyYrfbwPIO2s5KfQH2peGfnqiFNckVpUkVQQPYB
tmxSftrjx8bFkPH+U4wtXKXpvwY2A27AwZMT+KK9qiUbOp2r+5U7otErqw2GAFDd
NYq9N3tD6Mks8MAxWMkEvgFz0TgA/fKPMu8p9drkYOOn9VKv0ALBJcjfSh8S0J9M
mbWF2XDSDy7Qev72z9gMhGa4rM/06Wb+a1FGgLnQXiPKOlNPNY+0B7eY+UGoO/9u
SiZEN5y7JCTISb8BJsjbbWLLrr7TYQDvlGbHV07gc0x6eCB4K3xec3ZPfE6LCCMB
sPsfCBRTAgykrfYUTDXdSeZOu/sPF5Ln+PAonKls5Vk3De72uTG2U1gETZQv1AsU
GJJnBMf4XvReEQV5b3bE3FN6CTN6AWul3iFN/Z1tVOT2DnVvwpZ6wvAQzbV3flhz
rAW+8Qr6TJQwioXUUpApEkDwTlSY05zNMxuf5R1aJ4LDhXfXKhl5SNLwI558fGzi
GwDC0Gcbke9fqk601yEag4jpdlvJeDQiT4GPeBAu4QBLFtQUt27ax31d+iqWujbh
Jho9OYrh7QfBAfx1pvQrTRrKBr7rtOeXAHkkTELquYV8WX3Jo2abE413bwAFcmn1
fC4/9rdI/WasNupeYnv8ML9t57zQ4WAlS7zWsZF5bSSbEhE1vQS1UUSPV/kJ2jCI
gYpDUrMj//BRWhB7AIB/48ViQlHv4qfz3vx1QnG8EsrioIqy2saQKigfl5f9TwKR
6J6Mo0a5W5dc5RQ6XgDJT4aNI4DH7Kuix7qBxPdDTooM7DSo+arKpxxuCQub7GYS
1aV+8uSdI6PigL+v5Kxwe538uV8noUwaDWB8vmLK8Z0SPrPU1DjhoHfG+GOXbX2Q
thq88d0wl7UWl9dbqWsmsXzVhBUmzrYLKWwKga+1dTzCTncKnCgX40nfnLBqnFWc
SRpibhtJtfZudRQdB3WCQnAelJ257nKzmzKpGqW8UUqkcnQEjA605wVl1pe8m3qL
ECJY92MEaZvTeP2tEskCVIE1Bi1vsTS8wCLJAyv+C0jJ8npgzCkPjqGNVygvxAG9
Z/iUiRW1DcNz4NjWIbgw/EKgPJ9fnsqflcmZ8PYUDyEQvnqojXSarwqRuRSgMQro
2mPAO7vJtgEeilqV8vKz4VQ1ieUkvrh1ItuxtCHEAryhKWkC6xPOucFxjjbZ66P9
VIR5lVuZUTnhn2l5NRnIZ8rK3FC2Q3hluWMIe0ppNeuy3AYdTEUT+TwgLcrFMRj/
tCgfW8lsvlDnhGUKb3+d0NcyOQTXehXSvtVeF7l9jPMEqCiXJp7pVJimsfJOb6dU
zmzP1avsSOvEVw7ydHbn8Y+4BT6Qo20aY86jLUZzrK7UeEcFg7no86nvXGlGhnka
4Gpqp53R9///cRIur9V9XZewCh+ELZrDp8jVAV0B8ST4HZR/Qir18CkXUeSYfiZN
ZKgikWrNMH0DLjVPouTnI2Oiqx6MPnr9YS93hAQ6MNmJEXklTwDhWcbIVe+/fQf2
9T5oYa8TpLPkNGqCHXqujoN4idjweldyCy9oTQyeNhFHiO41ltBV2bCoP01m865G
AFBRkQxDxL0MEsLD0tVPWqIzLRaYXBVHZQxI0Pi3xgWGpqmKDjSfTADtwQIvtlop
G7T+IEgZH6i+7yvI7t0nTzuGIFRzkCrj7hRKw+D+kKjTedcXmFs5278fBxEvcvBh
nkzbIF+7kW1D7iRz3qRcF4jrH8XG+RWgFKcyKF5di40wk2Hrv2ld9a+jvnGkn1Rj
bQ/+M5UE3fB21Lb98wOyA6DQ0SdQBlE9R/YOKBDRffJ31hVN1Z3K3t+rhMtX+QP5
EVo0k4Ox7xyylAwsRTfouKoJX/3O3kmqDqwL42OW46p82a3lQJjsuV+JintaN05P
pKjyH3i80hYXg2x/iDdfNr9y7n1buChV+kpIRx4V3lJ1Bocq8+2DStlhVo1UutwV
3/vWTiTTyZjPTby9FLwJTRW1Azaj/bPkP/Ns/hGuiS0kr6L4ZowBZl075YLOj7hn
WY/fDwxw0BwBboKr6R4BNyMKwFxEEE7zqjTifvzHAumm/8rXFWhkjzrUSk4D+czn
DSAX3QPWKnLEC6bI2qN2IRQwReUzBQ7Zb+rhCDFqq5LguCwHf7OIX5P9eoxN7Px8
2GwGZUpCi4LOjLLbvMQKJKAYh/weLv2FqMTDNAolkEOZcw3JdZg3+2frpsY5Bir8
ZgBBubitzB9pcvBh8FK2YAIT6sWUKj0ujBCc+bBTaGfQQ/YrmBI2Oh88X+gXtUHU
kH6xRt0EoSbiBpg7fqdlu+TF2j0sFRRtNcjqd9rmqT2tZFjCO8lHIsDKs88WWVQA
mCHX/Ld4eVtXaEXrlW0jsXeeO7VhzlA1XBkOfpZUS1aPneJlL3B0kEx8QvnD1Vlg
boC8MaY6PSoaUCMAiNN1Wa5rRuq6uwbbzcr3OPUwbUEtT647VzUBNqY9g+dLPVdi
v+wRQ2mjbyrZpo2J3f4Ds3AtMEdhBg7IOtiAkOGSUW2fDsD7xU9HTUUNu4nuaTkM
imO/909fFQnc0rdMux3QmqPtD+q0wZK2ES7dvmaO8ZztMlGO8NPNWuDAyYAHuLLG
tRdUtIVXul9+VI2BBo+Z0RYOYYj7dFr8BMIsECGvM3vkcDRZtII/fmiAhFpZERQi
cpu9toGqJXPBhzo2475xih+CuQYqIJDQbA0+i9syvCcw1wCJqJrdT9omjRb5C8nR
AtQ0rcP+Kg1Q8+3wJBBcFiKBlPjG2t3Fv3BHNL0tcb3Y9PksnGh9d5irZmnmDt3A
7VB+3LidWslE9YXmRAjimZBiZc5DKe+nDm7G2uA4QuOeTYYvjDcO3SKJuCVdEhWk
3IjgybFEKiEfoKEPTlhLOshIil0H9c4E+rpqJrjcZ5Q4TougBk0Pnxpb7hZcNAuh
EWs32OZUH39L7Hga4nDAADkRVPMLdttXfspIUXIIaJhHpnR/sphXEGsRPdkTA9VS
e1KV9ydmJApmqyuAiJgcxHBkH1mADS3QJOIz/lzzYkPEZPMSg1s89yFAnd5VWYez
unCilEH+bkz2L8cqnKp9ej42vpL/cLmkvWWJqcLuA/P8SslWQfegbLCbF/T/BixW
YIzOqFDC/dNYLUtomU49V6GdEpFLZmjIn+0mwGlIguqy0SAwgXV4yCLjWWGRhK6Z
LNVgrUJQEnLZeYfEzXeHBHegGWV854E15aYycCUMiE0+V+40TAWXhrSZYl2RZ2nu
NuEkNJDYJbRhXHr9B3jEvCulfAOAZ8040IfwtibKoVYB8xhleYhw9BjkhV5AtqX4
9/3GNfCTb6oYoHNZgQRUjevGDo3KwDmNYcfPkukXDM3lU8tzSmgZp7GAN38m1zqo
6vpgeD/lYcGQEl3R5Cdm4hE6pDmVUgaWz6F0+KGv284d+UXGww1Io2zoUzE2DFK+
ZHDjt9Z2BSDseEm/YOaqjSkmsHAYti69oabrjOY6gVtNVHrFoOxJBpQteU6yyvnX
o+UaScTJ3UZuiH7r5xnBidwULxuIxSRr94nk1BXN+zMXsx9X3nkYt1UKV45B6dtC
AmWbJ3BuYhZXlqcTleINJjEWL91iC1suO0DIebiCtdSZ34Tg3W7g1zefBfL2YGUr
qRAlz2BRUNxoamEwW/Ycvij5GGgG/NxM37JMV/vJrf4+4b/c8EqkPDaVS8ro9Nz8
BSnur6KDblX+t8Bpbm3HLmyQg3PhC7oOKMsoxq0Ufi5cP2qqbCndClTLgFyifKiE
KcxmZyLg5cE7Mgu8NQ3QTawq2wPnEiZpigd5YvGR5JRr1668pdEqO2aOCeI+p7+L
lN/qVnc6xVLJ1wdGWrUJqnVi/4TbLXDKUYJmtxWFabMwVus5aIe8BLy794KrPvER
PhlqXCN0sgOnsq/Yk5DoBd6ZK9hnpaABpcd9OzdiHJMhvAG2dCV4M/TcXfYDnwFA
s+BhwPhqcOwuT1TFxek4UIoE6Pcssfg0KTTGaPi+52tZAx9DMGihH2SvB+ukMkPV
xgZyAmRPg7qDYVmaGyekWFAgozGp2caOZ/U4Nj/1+OMDTcZ1hXRWYxaB+pIcun05
LdvIodNh7UmGYutCMzmsRek2rMfZ6hAeVGQoNa2qGAnstPxG1mq6Xdcmi6r4sBQB
mtbQJnwez4rVI61QUCGYplo8pr/g0VF+w5AgF3K6o5xjLmCFGAfQgFVHRuwudYKC
6w3gYSrIYbnepC0kvR61pNtPtgotezP54tnY15V0emgTNQA2H+ORTWG7nlef4smT
f74f3w5q479VlD+Zj6m77guM25Az9BTug4U0Fj6qIjTL2IiFckTC9GBCQNNCJ6QA
VatdM2i/ybgWJfSTWw1vOAl4hXZKP3JVvuovf2ZQ/RyzGMWjmElrbNGgY6y+lC3U
WKMygw0fH9Gc5ITBwjZmK6MeFJnf/7MeqgrdjpXpHWx+x0nYsvd7JprmUOCO5pGH
LjepHDPts1Fc2jDzeKhHGupfS6tI9oJ+DLpTwih2qrY5uJnnh5hRiePgwD9k5ldP
nOifJOyPBazY+bK0psrId1VwEeTJ+WO+PnF8HTSiUG7EDI42oYnMpEnxvaGrcBmc
uwloLyB89nTsiya3lwFSuM1OwAI1YAAPDKas5cCiHcgeTKLOJGREZUEOPi14t6jl
35hku+UwzYQQ4BrbiWLjZSY4ctnmdymcFL/CulFb5N97Ok0WsVgy5AFRZ5A68rjK
fyxmfLJhMYKRF7a7XjOZooe5qmXKwxqZ12oUlj5R5TlO5sYsZVXX++HgVXneu4+V
tElc5jEVXBph6wvwuTgIoKnW5lr2zxFX+uJKvcx7pUEYFBNLmEqOvs2SqM37LlTF
UZtfnGX7ctLKVt1Ykf05H5O66K5in1LSwBegvRpaBp538OAK2cT6ePJkCEXNLXjk
1l2FfQMCNA5BZcH6UTffWGPK8OcvTayuFr9Hof0hTpnS/nJBfamxQ8WsnsWWgqG+
Yxr/2G0yp13b26PvMYg7qoymiUwfxuv39fLcdGkOlMl1GdnFSpRG85+fjdaAQn57
R18gGDY3qc7DHZFEaqVLRmNazvknNPfHXyrwxr1jwgXx2VZPi3U/CIsQdcUNb5fN
sd6htV0ed2BokYM+7a7DFMGUnVEgeq2IOYUtXR1dOiyJRMfYPNMIff6Bsx7B13hw
jeqUmiynU9TlBJy9XmraWBDBtwVN1KPndlJ84Hba9uAmmLiixwOuiEaAr0GauXDi
+2XySVUApfr9Z1Beh8kt2c9z9/4sdSgy5Vh5xRrrC6ErqPfkkkAATRlh5usFvPhe
PuNY4IczzVPhvjMfTjV62UKcR0wttoLMW/7RgR8gHysxahJlUdhykrN/WjiTElwa
x1Afh9YD/cgw84gt/De+IJU38bK/NvD9kY5MGZztkO0evqtah7cFeXxHxO1vmPRn
4WTlUbk3BguhR1hSoBGCKGXHNxqUhvZdLq5ePYlo0zxRZHIMm9GA+7NsxtbAd8oD
gqV2QEbuug9qNo5dP3gpAWPDE0NQy+sKGLpZ/+siOvMN34vhB3wzztsh/oSROnfN
OQdzFA71CDHLwxoqetz1KSbN00xNi/saeFLvzlVC8ixT7wvfbuAh69Cy+m0vZjDu
mc8Fvmssc9UucWtu/IjvwVq1ReeN562oTTPQMD98txC6AHwfrBzcJ0wIJHsg2hn+
ZSePpZJZqKDF22sOqd0ruZrD05JgfpUf4Sl3kz4d6d0moCmDEdBAnj7rw+YExDFQ
T+1sOtiTTUyAWCgqx6qn4wAMRibR0fek7MqqdrjaLxBl2zsekXk6ucPrBqoT/G9r
WSBSDCpH0i4DogMdrieRasrJ6+NXTFReEy1rScCNdB8oMveicp0A7n6vVPIOpRbO
oeADmcF8QDNPX06bRF5UbHKDse437gPQPMpgqVoOxZhp3BnhLQcAuZx/a9Bf26Dy
PXVgGLj6u5unXfmcDUeOxEk6qSC4BvhTuICHihHzFCEFSjpa7E/akf8yblGVo/+8
0xYVs3C/tjOYw4j+IV6ZcjfpxUub3uvXsjWOdLkj+h3dxwfe638jEPLW5YFbznS/
g7GuL0kXwHF05589DDdec8pGNfrNrst4tQMsrwyk1iXdjU/ZF4vDaim9gp3Xi35Z
kOTIk3Hy+su7ImseBr1P+CigP/ZxNIxEU1F3HKdjQ+YBHIFOJ3iUh7Z2BdqxWxv/
G+XSaElt5pQZxRVT3+Dmd6by6/jEmn3GfAcj6EdCaplVoJ2VrwxEoZYdxdkJ8zG9
H14wvQQVv9gXTMK/mp+SwsldahyINcR3pToa1y16aKPqc0neigDKFL23op7uhNyw
pwnCelzYwi7AnSoH1SZjYbS9cGLGI8w/+yXZmH18boweFf2tHZcyo+4bzWe8cxf+
Vugt+Px3gNtPHSAJA0xHj+xq7NCJ8G1Q2p+XnLAI2DP6hnbhuRFlObiooDw1TKSB
qkqXcgB/JN1F7N+P8eI7Xj3KXKkINnFuD25IEehxzaP+qZHPDnEUf1dh+P4CG+jd
jO59EJ9CezAIEGv/AYNN451YmUZt0K8Kjm6pL4J0zQweAQmgapTyn73C+pDplyxa
E8+7ypPLlfhqm/i4/7YhyxYkNCYralT5OR0bAj0DtAD30a3TyjeCHmiMBvhxAnC9
ufoQmr+hqIF0gnCZAmkugwczROOiHRbzEs8rpDYdc5Q=
`pragma protect end_protected

`endif // `ifndef _VF_AXI_SLV_SV_


