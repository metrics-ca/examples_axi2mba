//----------------------------------------------------------------------
/**
 * @file vf_mba_typed.sv
 * @brief Defines VF MBA typed class.
 */
/*
 * Copyright (C) 2009-2016 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_MBA_TYPED_SV_
`define _VF_MBA_TYPED_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
OSvAwSIi4/4A0S8+y98e4pbrRLnFhSWp+LB/93g+zZyATAvdYY6kHh9YZrQB9vAF
7IxLlH2xygf3P6YZspUgm+EADRTcCPyAFy2EYLwsOrxKdcTwraWhsvQGgjgAJ8Qh
NHu7wKYgVYxuBqycbTLgs1wykTdAzqXhovcdq9bM8waUPSPupKDeLp2WIXqpTR+5
ZHMnqTOqzlMmLny1SAJH1Z7GwXrVSsNs8HYg3ppnBtHYOq52839tI8BhZIcaMUY+
HV+MR5DeO09FShwnc38iImeHt/UqeGJf/jwOKMZHoigsN72noNZyF14yZN3OfIf6
UFGqyfEB3jWXjyKSNM2XKw==
`pragma protect data_block
+U3uIYRVKJ0gA2sddYhP+5erRAhoGEy9Gy2J/UtUSKM/Z9NDkk22ZbPRjkNkHEsJ
hHIhPWCys8paAPFXxmgOb+ktMjPr3z90YeOG9q8f1Y4oybSlZd1iA53H5EcfqGNf
dgsbeotEyAeQrrE2APsUEM233N3sKgwcBorOZdSnVV0exYcobUWCH6dlpKVPzuw3
s45lP5oY6iiHttopwiVzA5avN/a2CwYRFN9K0etYAAp492cGkO7hR08GG1U2X3eQ
j2HHAe0PBS/yvLSecx+JsCBt7smGLVs4mRoGu1OvDi4K9MOTD7A5MBcE7+9iGSCw
ptIiXVwHN75WvLM5hd0dphFj/dSFPcps5+PisIhaUQmW/fkKWaudY2QAvewy4aha
k7rwjZ4nkgOSqZCUzXhhUFAFFfvRy4/oQTezCvY2z0EL9fUQKWsHngqqQdbDBafk
hEgd/M6iCbf0MdTPRH4IT8akRO2Mp6XvgzR8Sf5FbtK8IwbptjdbCOVGxOCX0/7G
wQo/2XMKUXgTQnHIvTs64+yhw44dtMYlBZ5pvyNvlItHZSlkG6+FjPbPGA45wunR
6jrB9n7lY8kMVVE4YTgVldpIw5yJzNWmjPQ25EqvUk5DxH1A7lBpyLUQW1dLzRky
jA8pQuLIV1cHvNXCKB79C7ovJZ8TD0UjYkIx0ssz8dCISaObDRuccwnPnucoEdHm
9Xk8/D+HA+cRVRy17YX/dJEvp3ObVSW2ZxqZb5kJmqf4nJ/l0mPtgSVaHFKd7Mmo
qMUvcyS8fqcgmOQuXP1d5yBNOsAZjy90iZkyVWFA4Rd9YaUkaGJBk3fD/T3KsYfo
+jQvZZ+mqB46FX8nc6oQ5XUY0euKUnSI10nLxisiF5nuVkoGKqybGA5W5Oa2QdZR
duXGC20uu2BAXQT3EZp+xq13d+/PRCupU+KhEPQ65d1qNayOc+Uxns7XxPHv8QS+
K+nWlDkbtQ5PGNti4PUfADwbEqzJ2eqrXcgEDpoOsQN3/2WhXqtBjQRGsakImCwP
tfd07dsbrnfxoHA4j5iy2mw7BdfUEQEHqGl9hlTSCQdov0lz998PlviCIPaIsx8c
lVAMDedEeXzyyEFUCoI+Ig==
`pragma protect end_protected

`endif // `ifndef _VF_MBA_TYPED_SV_


