//----------------------------------------------------------------------
/**
 * @file vf_mba_sb_func.sv
 * @brief Defines VF MBA scoreboard access function class.
 */
/*
 * Copyright (C) 2007-2016 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VF_MBA_SB_FUNC_SV_
`define _VF_MBA_SB_FUNC_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
kWfpuwqK0ddI3XtIACKVgjXQpGJFojpcItm1pp/CXcWZcvByLiwMcJjNiFFPFGWG
sEGZIZFYLnZpZtHvAMqu/r17Fyim46OPfDtYRiASyg9HgURv8C3OzY7bPENQVdy8
DnAtWUbaTX15AJzIyD5Vr7Jc/NeLUPLVoj12aoTADWNgDyeaSA4DjAOT4rpb/EFk
hNEIqtPPjOmKtseVYevExmO07N8NjNdptLD4Og/N/F2ApirOl6sVR8dHjKHRY4D3
lu6gDnw4nY/bhMUqcEPy2USz1POEKyqHct5Py/9Gz7nxOKbAmkuwZroRXT6zF9uD
1Kj/8Y6Fkc0cjMBngdeCrw==
`pragma protect data_block
E4zpKz0WAISnQ3Q9HTKNtMeXweeAHmj2+Itw2k7hFK9XP5xsMeFmpOWJawfGoSGf
RJQYQmWCIGc7izc6E1k9X0dnl04NfGxRJmcZOrWDwuNxKRdRCsK1NCnVcWpUoyeP
G3OCwz7tAKyDgL1ARtRTZly5a7JXL1crQoqpXM/WroHi4R7YhF6873ccrFVMLIm4
9Zcyg0PDEgxEI9fLTDoLqzH350znLDgvscMH+rsIs7AU4T16cceRINSHP/qV9e8w
O3hTGBdbcJhuR8MByYmCOg4IklkfwSsrJsBEwCgfG6wgNFLAuq6rkK1Ovd+D4aQL
6RC3icy2A2awODMixsB8jHBZpUvQu4xcG1BX4zU8Pr3xMUxXUJKF03b9L8iA4wsJ
hdvlG/L0HiPiS9PMt0i26gyq2dY6Xe67bAy20X/mSCqThdUCkAJnuptwbWNDjS1L
rIbJGWmgxgZTIqQttiJAnUb6tBTzbDE8AobRhC0nD7Ge8IPXvVNKY813pMEUDgk0
LuvpW2DQ1gVfSQe4JTcm+fXJfd63q0rxZIoMTZbuODDNJFeC4DWT7x3jNKp/2/Ty
mWVzkTyudHlQpH9+P/ShyBVyKgrrr5xGm1HrxjcQeMMmx4kR+1+egQEYS4CjlrYW
RfGJbispLicNEAwn2/dp9p4QrsddaIA5ekYoP8//+2hUvm/ZcK4ZloT+xpagPvoy
ki1MG2ulKWPi3Z4Pi06o3Pjb0F0n6WG6zG22lQBs3sZMFW1VKoADuP6+A/kWFJW2
HarB9JNPPR72dKn5HqeEArF1wh/6PhEvkF4WzuNNXSu1yQL+7tFj2ARul0rDDNKz
Id9DTDygB5FQbyvF54B2rELcn/Mt1GNJhcIuGb20wzH91XhmLQUy2Oi3AoiWmJyX
LvCeqTUa03KVo2ly4J3Zkc0U05LZkH0oTAjo2MCQ1mSZrj8GUMqVAp8mk2JI5fji
vmI7rFLmKWwRB9B6umUErRrxDP1eFSMm+UWB+9LwAFLsJCw+TOExQOxTajlF68Ba
psUZtcr3RIX3C48tmLaYe2xBZ0HMUvXfbmegz260enpgCCoknvfjLjaTvmbjqT0l
tqYG2JFfhKFIGO/Autd+nKtzfkK3pCKdMKkBlnRPOVcC/4H+0h7lqVsHTzoK5Fl1
f+tPhfli5iYAUqvwwtclUSW6IZ5P3zKiJOYPbFE48h6/7ZrIaCpywg1S8sXKEIyt
eghzJEKl1dxgSGqpk1XdK/mQoTtnGv9D1je+aJBStXjO50HR54ZjXhsgfx7uZARS
6FN3217/CojoSehDPEEiahVQO2zeEN78THP1IhMv9TnrMwDOqV5sG7Y2oXV6zk8t
N0DDsesbP7JLv9kflRnN00duwSFmcc5kgJdYDhGNNg/crhr9LuPMuySUeo8My16k
TrKQW5rwNDN35ubSIcLLuvGiMe4QXQMUA7KVY5zaCJ1iNpMnk85lHBWDSGgHgCRW
i1BJhYmPUkQnyJm87OwEzHRfOD1qu6/43G0lLFIB9faf4unCf+OFL4rfkX+hurjs
urxH7wkONqkp/y1WeLFkjNIdENHiaRSAmZT1zetwHHDSGnMCj/dGbGWwWG8zt65O
+SB9ldyded7XwhxwcI6zMe57CxoVbC58N2yD8TDrcw9QEzdfpW7FHRtyG8nxvhmn
RrVgGDqAlQhsyq/+vr5ixH2xtxGWHgh1ezARHLQ5gy9cvuZ2ow12GDIxVfRODWdF
PrwgNYmNm/5tTEnXUssD9hN0DjHCg1iqwu8YJbC8jY+27bPzFNuiiTieTbfEDM2/
Q/EaS6XPVup54Xp/4MIOp3KeyxVqVO8oug/JFZlqGEAl/4V+iRi5F0vqjJ6LGHeU
Mi+IqoWpVXUHBoIa+7pk6Y2p83IEAkelUNmeafpPXj79NxClexnY4/k/J+5DFExc
4b6AFiiqqkX9IfKlw1RHhAC4IQUTMmMXPu+YMQ3U0YCI13r8XzVrGpSJGbumnydd
AdAFVECePfDIgIec+Qb/4OPxSrJIIIqMsVhucnG2ZNiloS/PB6Mudbdyty70diV+
8zfUIZgECPm7KTT9LgNQy5AtTG28JcFGYpk4EessCn+s92eQD7KJeYAL+BBFwQy+
CQhH7QDKpA49P1ToGhLlovq/xBiny/iTKICvue6J65wkmmuyLCBYnQ0Kr8LKjCeB
yLKd9igF6L78XQngbwE9VBrp216C9SgzBcdi4l0Zxjas1kaR8ALdPrIBT5lg0CQo
hHzW5CiGdiQZHajKnDJDWQL+X1GAqhR/4FaQ/DZSWKZZ/FqAN9QYr7hzTNwy1xdU
z2vSZYQT/wL3U8BPnKdu1X18N5fJyA629Vq2kF2j3vD+TAMT3nr62Y59+SL5fFEq
Fy49UIbTUsos8y3YpfBBpl7ib5LLzRqGmn6Pyj6lmdwhhvpaqJbpN4/zNi1GjHaE
NfNYmNLmuV67AGnwCiQ8OwxnH52O9EaWpLkM4X6hbEf5dta4kwGh5lnWbebbtKwy
s/VffICdhWHIGSBGIO5WHmWMjtI8nX37AxDuLjuK/oF6KaIAX+3SYKESsyCtzsTE
NhKpBE91LUJgB9C3UNl+DsrBpTe4qW92MC2OhX3P6FPQtJa2N3ypAeDO/i8ba81k
3yHoiUKo42nMqkwWYdG25KpYgHVWuyL9Imdvr7QGbOREggmlFBt7aAz93hF0AoAS
hyyKIGFFz+sfw4LeWz0ph96XqJnHodg+SKBJjce2LfgpZmZeZPbLjjxtHIAINgk+
kW3x7pengP3J4snQvVQ4FHO3h7qPXc3L3Et55DDa6nlz+AYy22duO4yn/4bnkyL5
XmUQRboxK57FHZjz2emhif9SkALEo1ZCmzKjIUCRmX3KzO9QdxgPMO/Oi47w5dvM
geYUToD2G8mPz4k/qZ7rqTMw58g2dyVkxJnRxX7wqgBo+2mJlWBaYB0RUB6rUiOA
skMFyQx3JH7D7domYuhQ4riX1hJXiCuglozVsMzOy38GuNjtN94JitoD1LIgrc8w
KnDStzBrT067BvNC6+Xzo3tDNaysCljHP+545+qCsEgs1ZdCCgTEcIKbsIL/byrm
mNTZBoiUlCHEStoWtf2+IVt9iyNAbLLJO1EBUBCXD1tGN27prZ2xlhHL2mwAT3Qv
kofvZmVSavpKgZDbiv0trxu7n9x+jr5GjjQ7as0cbYevpcXWVEAaRWJA+XWuBmuL
9UI2kwc42fe4nOA9B7ZbmUJqDV15rjT3O+gtzXwGONdbSmcek3VpAZ8jwh3GTusk
rr3xXgmDk/Dg/oqCTI8RhkgsR6iKwr55SAc3h5Lbya4MJkuTq7ETs2eIkHcBbwpe
hsaI/UjoEw2kSzjPj800QSR3+aDMTHqg0vRPvSgiuhziyCKHKuP7M/FE0oesAyJr
eO7SOxHTULF/k436CLst0mwCt/GLD3U1YZ12NDa6rov4iSOEWoLCxCwXvhf3cttW
x3Qonirizhf/xfecC9EpuY0LfMdgD++q7VAts0IOkuin6VOkBiqD0X8j5XDTjo8o
S5daWHNQ167AlzDsor//jk7pa9y8VhRr6mVB6Wrhel6iHF04AnY/9P/17lJFTguN
mbqryo7l9xnqc5919SzHYKnSUH+udEYrUGvcF0YGJQrNJJWRFQuLs3BauS+YMJla
22cubPWuPULdhm9JWVq1XkGomrrZBPEnVQ4EfXIiSnSRO49B9WPMdWwwmpzsiZwd
U75eSbhIrlwxe4ju+jo0N906/VpvFWaFTe8w6koeWcri5Ig5vlt44ZKeMzfhExT/
EAOUSUZVe7a0+0/jMMMxLvjPgWS0gy+9wbY+QMAc9yPAED66nM+8t/njfSgVPt81
YReG0h5IFXPWR2alf1z9qh11zuM/LkuFU6N3wsfUMQgVypimLY42zMxepw1Rv8pe
9g5aE3mpklB2fztyWvckU6BhQM9wL+GgD6IO3z5Xd3NtooQq8SImo/x/OUs2bAD3
zsac9TM/BvDgKqLd8RW9oKpV7x/DHKMwyI8jV7hhP2CSrejW9XPOdeHTdZzBm9o6
SmNH3evqgrgwnv9OO/N7zKIdT77r6meeqyfUJK8SOtgUBkkAyP5FhkHhlLfjv3lH
Z5uKnDDQS6vju4AWs2eT6eaHDBRwBhbAUdln5CBByJV3K2CzW3dhZs/vDjl/dKgA
RmhZo22iMRwZMUA56amEdzMofgzAKY6WQTnr5D/j/tWbf81Iv9btYmMsWQZETFjX
KqOa9zsO7LL26kMdNfMUb4I6WbMBz2h4q3x/e/zPq3fEI1HRR/fpxLRQmWdMy7GI
LwLAvRs2Juci//ofq+BfIMoN8QyQqlwC1BhoC+t8qrMAu1KZA/f43P6FQXGNKNIB
EYkkp8kL+Gm6MoylIVyo9x1/kum7ICOJx5tkHGQmUP4vuxUSmlYwqkafALgBl8N5
G+g8U3m7bjLuZJuPsYkybA42Zq6iYsDZmnVjRsl1/fndtNRcMqvZ+Ur946E2t8Pe
yv30Mqr1RF3HWfulTS4KcfZU+qtqpAd/zOKK1oq4tnjkjGnKbX4TfY5JsB6YKeIN
Nk9dsId4QtIu3L8AZIggsucbWd6DUToky4KANiMCifRFURJAuP+JstU42EbHMAO+
amS5yuempK+PpbSczZvFjhmptP+EGFISghTXEzMe6xsUyzUt6uSclyiPRiX0pTN1
4R1AdDyCoM2tihzbq8S9IuJeKM4LXI5rImIl/F0bqAi94Fgp4etD2AzRSkG2EEck
WkCuMgHg/88jaOW+BzYlXwVSIM/VKBtHvSxdkozPJe/Favx7r99x/aOUfhOnuOJT
GZZNS4jgi/UcPYp44Pds14qt/HxhVla1OvNPvstLCA0OLyF1Tfu9hd1w+ygDhwuC
4qmno0unlB7lM9H2KKNGEVNO8zYgK0puekcYkz2Mun5yHsKzZq7U8LLQ2RO243r7
yWwl2FV8H7Sc0Be59Q5kg/QYS1I0r/bfYMbWOrLiAZoWLjRp3xRvaSBNsi0YnYN6
m7YnePSIylpIvEooGqlozIYN24i1hoKW1LuFzDzec1nJHkkjpiGQDkp2COkjNoHc
QdoTxmQkfCYUfAZJ5IvMxOMiFcAjmTEvxQCXU3CfFyNtlKbxKRl7FPsy/VGLpMgh
cXaA4tQroCY/95oSDjd2fxZSDI2atF5wePUOZXTCc4LOAXmy2Y/+IUyRNoYOLWwn
VyXH1ds6BUfyUqlShYeuxr3BDdeOG+De0rL28DFOORGoNdNjBNYsXGijCMyn0icD
yxD1YwLpsoMDmCOPnIbTKA/p7xY+rhPHd/e9k8gr7cXhFIqwIicaYIBY9NVGtFkr
3muQy041TKDiFJqA1JrJMlNeXSLaB/eJ7me8ljAHksjqnjjplySezPZOTb0ucNC5
Kc9zYCOpYPTNAW42Owz7r8jVFqPqHhH4ok94nOmbgx0upCZi/83TKRuX8PepSMvf
Ln0Z457PU3pCbjoRwCfJuR6/lO76rwAJL/JVemw+6ODN9+yuXyVvdxzqSkCMSW7n
+a9k3UEKKBUdj89kL+Pt9KVWDM1TWLhOrqsU9fGojWbf5TkhcQ1l7g9xEYHLE65x
wmwWL5/0odcGAjeNoVBoBgC2tiYLyLw2r42dCqxTrrzbN01IPPEu1BVdt8W4DygM
ptSGF5V/W18bLR1bpTPvzqg+r+BtqQ05yl95QNoxfM2qg8Umjqg1ECHlIkv2xxAa
vetKzY7//qcaFpRhKQs9BXySOOgGbHMzN5+QCXqTHo/63VuOC7jCAlW8por4Ekrs
5bdpUfLqU2lIVJnlJugwtSvxK6N1KmzvHB4UNpCEmTZ/aCCx3pHzKmOJcuvZ8RRV
zRjCcD/S4ikZSXrw8jNZb+HNZVxdy6f8Zn3XoF99zN3+mq18TDSoaWs5a92uF/U0
sTO2hDNR2uNcJFG3bIA9tyIDRx96ZfWxwIFKUKhVl4ONb/2ulUVJgxfoFioXm/r2
+ntDN+vaSzd62nOQwPqw5mvPYWcXhsl5iWa5mUrTJgD+VRxBf9JjRYrGvhSz9vYr
TS98cu0wbkdbHdmuX3fNGqUx0oU7mvaMI4vwz/fylEAaCTXlaq4TeI75c+k/C9Lc
k/NdQ3B7U3QT/GgFBBhPoGHUGQe3zEXqxvX6UuEmXVPTeZsUx8Hx7DQxwuCkU6Tk
dMd9eZpc9eTP3TM0DsBABySlbJh6XNCkTSd1Rj3gyaFonGHv8DMIMJ+i2lEpuXib
uMFXTUeKsCkSaWINT5eW5cT3TKNDIk6cwLifrD9ZI/NfLxW8F8z5wI/LTLys0hVs
/MZ4fu2E/8K1fLlPgokrlLY3OyvEMq9GqjHzLComxxf8ELdnGSJAhM0fKqfwwA5R
9wg/FNaO8RvLlGvDZGmqrykMpWupBm6G0WnOQbHUSzgoOBrpTs38AdMx5Hu4l5HU
tvVVV8kHFu3qKz6YnubQHehpIjgFur/FAVfFD+8cVV+nSvSl1gSyEjr6IQvGPdLr
tzxIX5Y9G/1PnTPrm0NVd8vAE2lGHlgEV5dsOdcrXlew7If1trn02fnAdymuHjAv
dpm2xPABlwaPitxFGFXorK9aUTk3TVtaDCpPidmoRdyFQtCtAvS8S5569t7pHecO
wp8yzr+Gv7txmD3zqM7eKgXfGPtwfbjVNaRFFYYBb2zBAD7QUrGpw6sIEl48cTB4
oSbfpABVEKSFqqkgGNvqgyFYVGSRIgxK/J4BOjzJvEhY1pfELdqVTY+JeFkOxre6
dZrH6+bSm6rRHv5wHzvaLhDiFrhudM0XmPHg2wLQBM+5q2s4jxxWdtc/B2Vo6wPF
LjmbjIMXXl6v4V49GW8X5xg1T2Oll8u18NdmC8uiB9+ank7kV8/h5h7AKGwqumON
EUaYZnNPkYJBY6KjtuoHjhxdU5hxglPTfz/rsQci53gyH2VPciIWzdCqBKfYSS5V
eeqvnJFy78KDogRn0N95/VOA9oMZP24iH3InI2g8cY7CeNELX9rLmuLIdksr8Ep3
V3QQ4nN6L09liXAEX359QJdVtHoFcQfBFGoSMduisg3jo1H85Dh9AQKJ8YQHD0ze
2di6JL41PAoVbXbX17Isxl+i69krDu/9nct/OJvwTaLdgIUcUDaLFKY0CR0rCvyy
tS9o6DT9BG0V3cPi/MNjzK1P241dL1zjZ/fQ8GlePLqhjAYsANqzmO2M6UXjhjJE
kN0r5qMEb1T8Ji13s3sPD/RHbGzV//um7EqUJVnR6QNO49zzXxX5QQjrVd1XoBfA
aTawfQzbswqQOstC/hBwyLXW0bNjFVbzK4+5rNgDlfKIObtW3UVidZdlbH/FSb09
LoAJEaiPbQsQg/zvjv5u2aAP1VKf3gVrcySG+ZOxALGjsUecEAM94i4uoNBFMt5/
bN1XBnbkdwCDelm0J2i9bT6wMZECSJwNkaEVAzkAav1LMD8nkqlMgbginlLwl1vK
94jlBYTKRZ6/l6bUQJPgSvW+4+FqhgFYhyvCQ9XtGfgNwLqS1ZE1X3NJP1S+xU9+
cxW/J9XyfQfMhpBsohI8fWG2ZGGIFoT/dEGptTv2jnnOE4cNK7prYrBLlVGEczX4
2D4xEjHQ068hBercmEQdz1EdZE/17dU4i03Ry74oH8K3Snn698Hc4pK2mr7Obtq3
UFWmPZCxETivn9X6/YC4oz8SkXO/wiMA+TwLvYqmFyUFMFX2Pr+Kb1p16+tPmKtt
d7c2UyWKNEbUDcgOtxOlwTm3IBsRSMl0N3uFLmtwswZIZMoQa9UNvFYSbNP4gMlR
TrV2S/AiiRel1eKZr0w/S53ZIFJCsMTSKyaRwuCoNWt/Xlq1OyVIlqzLpijnT5sd
ojnDXbD3waKJPhkJw54Y0iiFI1zLPg7jgCRchljNsoVRsDO9rufE6HYnuVNU383L
qL6q0or1IA7qvwrgIGyoMPLH5CKzBJ0FReWVjkSnm1CEkQpC3l4WM9xQXUMlIZP+
vZj7tBD9CvF6UDf7sHKThz36FwURlfkJEOKXBWID60SS9aaw0jfoTMgfpturNoFs
jxCUcalk/xlbgl0RAXD5bjbWCPRG5vVv0xva9Bo4s3MliD2XVjyY1Dq/c4mSCLMV
5ij3lJQnsWUraH1Irjqsfn/Lfh5p8vZSa7yOvkBwAgCYZNIlTl5I13vnqOJuB69/
AjawOr6sCIAOh1h7s8TZ1a5SDw1o9tV4NKS6ZooF/Q8FHTUt+TmrHQmHTvNn5hNc
xC2Yn1QERCl021mS7pMI152xodqKX1IWpBi+bmsnFqh9VLK8XLsBBOId9Ki0NI3T
dNyJ3Zo9zuHJUV2FICc8TnMTMwXker8PKF63JuY7S4VHmW4jRLnfYYj9KBvmOEFA
nHkU7fCdVyU9rUymn7RYt4fWv26VXGu/a8fYI8q1sk0sMxBbaZiR3DhaUhWSzNrM
TxAZEwe2ZH6vmZNWax9gxgLRd5I/N60TFvrT/C9V6PyJ/0zO7VYvttZL4G5iBAfM
wTXqog50usbfFpTus0u0mIcx9Wp5jvQrOhS/+sPUN5elSdfHbGGF+QfQZi1OMIQS
IeI3BT5CQmoInmFChY7MC3vLbOX0ZhA0jbHz4Wj+f6t5FANuouSwtLmkaNdl2Ioo
Ye6EIORuYtjG2lNd9fE82xdyJG3gZL1rVndU9XBKah+Tb0wKy4nRV0CfvPNR70qz
wGhlGUBpLYgFRPEErXnfsM8wkyRkzZvJ+6FEhArbFtWw3MtI5xhWa2wxgswrPuXo
LX20go5yzfgBAgW5GEd/+qO+SVqAOUP1S8WzA3OIyhoeHRIX88QGkZtqV3CtJzeS
RQHtVj8B1fsN0/wc/g667E12EEbo67Cxt92YOn4H2EgC+ANq58Nj+QeDcqgyj8Mq
LOyqGwR+he/Kcu7GtyvYZOQqpU2Sgrp+ao1hcTsHKur6ImDGPF7WT350KcZTVfXn
xcbji7ZO0YqinadLpY2s8f+ZAAV+2Rb3eDaRX4DtE9XQpeinVJfNeF8uo0v2p6uw
U29/qFl61hEBydcArnkEG8xTMBZGzLusHOHSj3FhBonKT6xw0lzm5QOHE+uokC/e
1q4zS7tB0Z7tZJ6VTnzc0Av/pyzJFY2Smc1o1IxMCVKeW0lnyOHQE1GSGNsVlLqm
67WjaMQc2ZxKfD+Mrho53dkGHsCSyxFmDhHbDTyIv6w1AIOEvm1Mn9ldFtC/7/n5
VRMgHPVTMjg4DJs2LBSVE4t0TTk2WbQfnHDm+n16eqcZK/lzvOcx/FnEvdYx8jZ0
Tex35Z8jpLHTz+ns3/amdhGNyChgw4owjloRzaKXj6LceLC2wxH+t00kDqeF4dVK
3J5XsFadazRyUK0fVERYHLzkb6SgeA0E0LwRNfSNuN/OkjjFNNHm/+kyV+UtJzMe
E3Narw263BP3GqayziSDehZO9ydygaGRETE0uDeOj6us7TSkxi2o+zto+jGiHoSv
iInpx8vhQxhClsJKwrFBFDKbbnkVqz/dPrBdH9ncAjL3r1fd0gXGeTZ5odc+rU2w
7Zyvq+cQERkY7QhmYGs8/hGvjap0fixJvclirhJM8r1Gnrv/Zg1F0MObbDnm22nX
zAdayAOmGAr2zSltnBANAgVrjNEHt+jcLZ/veAkoK5UPgbomKAgllP24nYzcOn31
Zoq9R/hrAaQlA3lvJYq2bdtGFYGCdBahvXbOdfcGrkwCZfMb3xurD9cCmOryRg9B
w4nbgBpasghX3M5/wXC2ZwfaAaYYfEXBK5DoDNghdtaS6zS8PcaWT7IlVT8JKsn5
Ki3QxF6MuT/EA8olVSEziTsMBqLj8HaatK4dYsVRJDRigi1MoOdJj5XDFwZ18wfa
1PDiAwcn0LQ7Ar1kSo3FEVNfDGxfVup6TxcuHaCf+zKiUL6b/rrYCRtnItq33DaW
YwvluTtUtKlfORmx0nEuXJny2MMUHRFVrx/OpAqy2Uq9VaGpbsFXgNmQsN7ZjNlc
JEkHacMEpkZBi8JoZioLuEcMSkLaYYTB5WBMjn8WObdnuR+uNsbXEopTGXq6R1Nm
djGkJqbNK9YwiFI47ShSw7T+/BBAmCcz2lQLlbnT54MWMTnEC6MoyvKgImYo+mXQ
S5srD49EDwSGlPxtGipEU4aXHePNg5uV83mnMiXYhdVIOcxj6jH7qPC2eeczvjnU
wQz581gxEueoY+5jF5KcLR0jP8W7K0i6vtPu6NpCnSz6QF1TGwCHIOQUnv6iGSEx
nHlqvQqeo73CRxyve009+SrOG0v0BQnWEEDYFcGCjRKlE3jbQGRg3xvikU+RJ2p9
duBcFKqumGOCRN409OOSp/5MuR3YGSUl3K2JAUU+ejuM1waRWeahe0Xs9Gd7qxy8
YfT6jwJhs/eOStiQDmecUhVJ96AH5ORgu+0duYUzGemUrJWYcrTHga2D4BGnrUOF
YPeG59brhRGkZNW5WvI1wNdMj79G0O6yUymDGc+dbohtdywUoGmtGGJMyXPIVK/x
LEQgU5RM/5PrlFuvj4NPQvgW17/Sasm/wtuJGk9wywmq1mivOnuUt8u82dYA4oJV
o7ApCIDWgzdyOltVwEBfiH6s8jHek4lwJTjs5LWlaVFbM80Gigq8NQ2ivqGXpX4o
O/h7YbqCOY2gtVrcJrY+03cylsHaRKqpNNbK5FGQNR+z4WtjVZ7vutuau8XfdMzb
mN2+ig+Y/Ir88Sp5lHELuEDM6OM5eeBD3rFHSEiSC6pboLDen1MHkN9sQdy/BKBH
i8Ls3Gs+bCZXGmJafFWX4Al/Af8LH/N5g8bILFH+ParD/jKmihAS33LZXQ8XcwxG
UsNYlqN9hBfRHRAInuYQ4sU+HHQX+lA3vLKgncbhJsPmhJojc4Zka1zuSLsFIHEj
cusNcgRu+vQN8JtXF29qgg4G9MmEZj3rlzPPDYI5Z1tVIapv/SVfjadceL9q8IEH
ziE7oOhRq/OdlLtinUMW1PjCp+4xQq8TcMLcUUJ9LT1C3ZwK6Zxf5jH2CNmgGqui
QH6iWHDPkN/GlRg9C7D9xX0UnVLTKhP/3d6BacCyzLpopWBPtfw4SzUDOKBxnHR+
+O4k+fg2KHLffnePK7rjPYFgcPfa3ibCRhkxaIDejcJ7t34rIGNqtmreCKUrsua2
8iT5WbSGGXHzHbQfRoWQ7vrtPXS1HywVeMZNfKZGMoO7/DU7gLN8/hURJZw4j8lM
0Lu4yPACVXjAliquIzAIjTTYmwydsm7p5ExHmsDRf/ntDLArnrldJpSldrQUtFA4
DxX3obV2oRhK68Y3LS78o4NCnTGrKJ6Ff8w8/5VYfJESslkIBI36sdf6pmXA1D2b
QrnUxvOYzSMJmHRARynysCtAf9sBo+Fno5VrkF5J6uIG62co6k40L0q4sXSWoSQ0
WqLtUMXzpaJ+4CeZNrDr//xIHm+Msi+gZfzd1SMaRT/D8m6KXXb7LPHtqQZHvXc/
TX7ZGYorn1Z+1FOWLE8sEv20wFJshmBMrwL5CApMrBC+TEc2pVpaZgY4hlGuo+fl
XysShbXmVrcZWiyjO1U0ofmrlXmbpVyhaPpaFeG+nHQCE2SLgjDmbxr04Iu3/lLD
uXCjw9XNMRPdNuSFDBSMqX8+JHqq25xxdqu+ruc/Rq4McKpyLlgDv/Lr0WRa76a1
BQaGYDXYKb+POTdRjpEYxsb1DqMU487jv6CR1T5Dh+ulFAUHwg6i/LVogMeqWa/R
NJrFF1rjXKsC3LT0FlyMGY+KJEZyB2pjNed5T+j7IhwVtMYdf5vRfisq/0mByZfI
DrZ9X11pEztgZkSFmf/AaDR1vzq8k7R1nJQUXbZ2VcUPq2B6hnYoNcghipx2LTxQ
ODTCLCiBBsVph1ObC+L3n1nnJi8+iHtvU22sz8gYJri7KE3OAgmzD7bLf65xx4Ak
pM42C9LgbF/kclOZzyhwRIJdLTMYXj9Dek8yuklTblUxe2pLzIJ3RePrPKk0RC5I
VnDmb3UPYR6P95udGgLjfyItejS+8w392IBohImWisfkLli9nyju6u7OE1ZpqrJ/
jLoxHXbpLjHwUWo6r5D6SLHWIXHn+OZk+Qiczip5qFrwIHuJB+uk9eT3y3MgxF+2
ul1O9pOwiHjurWcCi0T4pr+3lSmqGqVD/Cc/kMvWkp4E3fdlG7WuzWBUXcUzjAdI
EoYKa6jTXV1mF3hzkzBMm+0LcL10IDGzm29a2s+i8azm59HmvXfQ9PjnjGPoMqlG
NvN98UPTLhB/J7IzeJsz4ZcxNhlknb1dCa3p3BGw3cFp77qI9Rz+uiBzBm4QR0jI
1aF166NGP1vxGAH5ZP2PRVte+biWBxaMttfENs70pJKZb8G3+458JOXyL2rjSeGr
S0NNQEtoenVCNZhu+zH+cJQcOtV4LlRqFTV7NvzG73B9UYHQ7fZ+DKnCdhget1zc
gJzJsJ/WQ0GAu8GYzGUliW7KYQB8BbLZN8fl3CNWowUgz20Rl1MjJTnPrhVWUazK
IwaCaFYLu/e8Mf+NX/uErDi4Kh/frImDyHplZmBItEu7Vrxcj0Nuc5jXMtBwpUdT
Jzfh/lme8dc8QxncMmNFgdPv01XKxX7oN3Q0p0WYxqm7LnCvCXtcpKAl6VuB9w8L
nd/aaypo16hGsCNmruLa2ODe434ResPAjgZjydZ5uGL+107BZv7WIMW+O6KuJcJe
wMxb+4CwiDuaj+NTnyV50HHGPQwGdYCrd6wPqgw8Qxec8LQD+sCN1C/8U8rUi/o/
mv0V9ZeLmvzPGraPzDqyZ51SZdaFZCDb4iR5W5fEsKuMq+x9ckvwU6FYH0CBUUBz
FTwonbhOVulrJryFguLf/6MTjYW1L3b5FU9q6sJpeonA+DuXhmFH04M3eGHNlvrS
H6sPMLhwhS9SeKGYS/lSPzuQf6YBGrR/ced4zwo2VAbSoNaBK4C3plNVkAiwl/St
H0O4XRdgZOscSvsLFEM52jcpBZ4idm1uAiiSDqo99AuSWjxmBoUpXvdDvUeOTVj/
u7UWCsY7Q6o/Ic6F5eePgBYt3W0oJtYgbjkP12F28n0=
`pragma protect end_protected

`endif // `ifndef _VF_MBA_SB_FUNC_SV_


