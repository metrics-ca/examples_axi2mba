//----------------------------------------------------------------------
/**
 * @file vflib.sv
 * @brief Defines SystemVerilog VF Library.
 */
/*
 * Copyright (C) 2009-2011 Verifore, Inc.
 * All rights reserved. Property of Verifore, Inc.
 * Restricted rights to use, duplicate or disclose
 * this code are granted through contract.
 */
//----------------------------------------------------------------------
`ifndef _VFLIB_SV_
`define _VFLIB_SV_
`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="dvlencrypt"
`pragma protect encrypt_agent_info="Metrics Design Automation Inc. P1735 encryptor tool"
`pragma protect author="author-a"
`pragma protect author_info="author-a-details"
`pragma protect data_method="aes256-cbc"
`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_keyname="DSim"
`pragma protect key_method="rsa"
`pragma protect key_block
gHmkj/lvlBtNcfIoK7Qo3ZtCx/nOxVYQCUzocLivF2A9TXoU5pYs3g8wbvyeDN1+
WhFV3+eBtjKUKEnq1eztR3u01QibmrkKF+DWK2D62wDQjNyDfPxA+xCGvtgWtlfc
hdET319PqWqGVUeOH/lG/r38mMHOOPKVmp7YFgERct5/gZOY7NcEs/Bc2b3q65qO
yhFFZE+YZw6DteW2bQA4bYNTs9rnlTsGytdtfSVMSRxe6TOPo8cblZwPLt1yhsDc
s2bvIOmEX3iRD7QbVBYmjyLIy8yVw6DbajMUnKWp6WOHz3csCi1QdnzdHf76AVyM
mKkZFquKFbReLUcHRydiLQ==
`pragma protect data_block
ksvsXd1c1OJ29si+h8uiTo+nTiDytYknPsiU+9gv+30J98EetVspcZCLWc+uf7g9
l9hh8tD+Z3haGfSzDn0K45/t/zz9/Y8Vo3BhmL/2F5W6bbwCX4iaAXaUc0DLoW+p
A0S5Sa8DG8UpobmFmKSRnMpKJHAuRfG0+NVouK4NtFvOA2QEyPU415uaO6y332Zc
tDXNmEtMTVuqgCkmoEbPz0VlkhBmqSXP79A3D9ftAyyCqG0L57GPqqFyBIX3uFHY
XM8B9cdWYEjvDZvvN0CzXp947bged4uJYJ2O4yemKbOx+nqz872vZo6IjzDxHs9d
sKJODiW592pytQm0+8iK+3b2XUNslUTcifV0DCnNm2Sb0EFbcIJ8HFutlJsdr5Dn
0UpRYoIarpsBf5tzj4PwyBsFnJ03QXedGSaIsD0Bo5wKaUb8GeVzmcV9OOrVUECA
S0i2QOKb0lKs459zEAz6V/EjmvWAZk+bY1lmOybPdqR4I7ZiNQjX4QmXL/A0q2QG
GFfYBX+6dsC73YMV99yxuXpkyGeDghY9AAyu/t9R3G9A2k9Udi2lC3oYzHuw0cWi
ZRNKEATe3dJhVZE/aqsUGQ7OHlXslwf1VncoMbJBdix1Nv/Lo/iK8+3OuMvUeEyW
rlBmRFQYlS9zldCRadxPNV6D4BpT0sMKUSoD426+xwnsHHQDndPxjdqYTcAp0abG
9oec2BAw4pRll8yOMIb6qqJnfY3rR+6/PShQ35TPxkXmr6mmisDBfbFSMvvkd7oH
7ddnIkaofUc/M7RlC21mY93XVPd8gTJzziM7uJt9BGU7Jfwawqtf3zOGrPqL/O8e
ktB7kZc070cxIp9/jHqNgO8H3/4fF+YsLRjUw/vfo24R/MKvCT/mVEGRTEpuK33V
7TxYvZk8nwBiO5a8KxPyvClnz7cVyjcH2tkEUVkrv2JqGdfMU7lH8bjKatCweLSJ
iNqZTCBB4ppjOWfLH1FvNLHRo+TeW82Vf+BQdNFVJWvwhHpybPhD9tsLLSXpT++R
xaLbpWdbLDvGl/yQiHSXWgJjJQpRaC3U3e4E3daP4IkZ+LQVEB//BsU17QXLdaAs
4P2XtVSPW17qNu5oC5RnZ2snMJxuCSxq6EKRhFsUbwbI8JeGsxcMq9FH8ZxFdohC
+fd06tYjr8tVBG7vpRS5k4fHJD+dwf7dPBzP9QteQ/7sEuB0j7byj6CsQxvGRcfl
2d1NelB3Cy1qn5gwfnNqmZCuWQwRQnW/Oh1r2gvhN93TBdaxTCoXL91Kd7RHGhx4
0f1IKre1oaiS9x+XrcuZTrSL+akCbzoH/njqElJ5Jb5zSLj+UgJnfzLEh4ZXqaoU
KWxYRxqb3AyFhsXNJaC52XZMJBMb7kijeLrGx8V4Xi+7wxaMHSe9L6PmfMM2PUKA
+8YZAXe829FqcmNkmdBw1xn3iDUUHwqeml7LgPUjqFuXErujvFC5Tpm0i1tSHoce
HSAcSZA0QVN/ojx9gMWu++hqz70L0gylBG5auPWgbnaRxcL3la25Ai4ulJ9a8AJ5
jHOtjFrBhMf5K6UobfWUYIFMznz1mrrj17vHMnYzl6fv2l/mHJIdrc/7MUrrgP+P
z6/hJq+zhMbVgvYYraPP1PrqG7/D/2wEaGeBCLMEPy9bw4gbCdWkFVDaCIjeod4a
qqBF/ZojDJtCbXy4zoAloaVz36pO/BH3rpzsqpQDIxBEUNNTQplv9qQWmRdiLCo6
nLcqH1TYvEr1JM0OE72GeAWubBajeI2wGV1fTh1K5nnbEJgRVNfcAhzShADHvrDU
/Zugs00fcGwHGLsuvhdgqY8w+5oYVZDA494nceR5X4xBOtsnhGlYwV7pZKsu5aCC
/vRxhsTY2J5S1XnIMG3DUbfkyAyeb4uzMotzOYY6KB+s+XuA0ptpRlDAs3InCW+P
j2/Lu+syRmynyGQLHvr4YHyme3y0/X/++BaISf8c9ejHxyMpsLSHIi/IPeZmBuht
vPnay/myHSyqN0kES0ND7TjStpZDL7PqVxqMkcSaXLSEaLMRlhMczYXP9YDuqsz0
hg52Ey11C3jpaSgF15C/hi5MELnO7w8mOzyvChVqeej5bScBvLVc407MwAUPmqy9
/HKeDGzjBjX9PYg8nhvx91Tg9a3wpKCTI5DCkfg6L87ME6OpspWn845w5IWVJxrb
zkukGb/9xUSc10VL4cHqI1sB+i/ORhWpoW7qhT67ijw4Nwx+cJRFqP6chp4/U6xW
IZgJB4hbRD848HOzt/Jg7jxgMhXaHUrskA9AHqJG+w3nZNnFRtCr2sYWBM3mzjvP
72JUfQ9K4eEY0mpUOL92Oz4uL5nEBZpxRGU3x2O2TY/JjXnLJbk3mxDtt49OTSW9
njQgGOkTVtQJLew93PI3RG9hWjuaKglt2w/k+yFb0s0bigi1/9OywPEWs7eJSBRW
ISFaNC2SQnwhcy0RD3pVmJK2GOMI9J2EQ6mz7BbT2dNX/Kgbs4diPZo/EisAVitH
XioFNdnTdAckhG76GBUrSxSExrBHAOs5cSk2V+4BuqjEhhY7W7dms5R2f7J9R7/0
zIAqmiYK1Y8ajZW2WwayzpXRnH2GpKBcsFtQNc+lcJYjxz4tJqwdLv7tsSEd5xyw
iE+jf091Xcd+fpJ/xO9VJjMUKDUQ1QcieQM8xYacnQJMbY5freK+biJLC9ODmTVG
SHOUtseQeGHMujskYZp9IMskaSzGgxWdDsuDS48d2zwNPe092AeRS5eQ48hvA2cG
Smfi7afbgVfpIPsU5sBl/mr8Ps5UQeqy71zx3OzH3Bo9IIlGYZeULsZ2cUDySrJw
AU52JkguBNLfXufaV12ajfb5ZhNIn1O1ITuf3KqHA7TEKACzdDwoBMoNQSQiVOg6
LZZO+GaPPoSDZFbbOfE/EBLZkXBDEFY2LCMVM1mFoUvPUNXP+UxV7KmumxqCb0p1
t4CV2tXn29uZyGDb4JWFWKXgPW8Qde2tinroI+wO3fzfMZGGZE642K3STCG3wq1g
U6XRESxg9cMroQxuqHS+RX9itlQaol8e5DL74nq9UNSDoi+N/2vHpMXyaHsexHqJ
fs2ea4E3sr/pR4wxRyejBC2WT4zQB+T8Mg1uUv10uRe7kW+z/XJWsJjCEObZYCXn
s31Q6Z6kxsXg15i5AYZk6vvI2P11OSmwXBbSwMZVzcUqf73RHwRN9IuI8/PlN03n
t/TypQL7HQ2SnGtDRbA2BB/wkgDa5erROF9k5WThcPJvn5FJgLDTWSsM9FfesD+f
XbhDFa2T6TiXYIDIjftQGUMHnRjSbdXhPP/IXeUb2flRESSBkouTDjOkPt1sUXQO
9/x8HZC8RCZmVmpFPz0nzANLVGSRUjPltUvxQE5S1ebd/6BcLbxI5jIKRRv3LXHa
5dqZZ63HlQgXOwVtspAG9jQnmfGH3kTPpxcoKND39G9aMCWXcx3j97LRnurw3T6e
Yej3mXBNfp8NIXpFdZTipXUyAcfA8ZfqN9MvIXcJILFRQJQKfvZHDzoNlOliJI1B
DaOzxocIYhF/HCE3ATEXaeAezyJXqENyNLyP2GHfEGmZEwd2ixu7fmM9qLZCeWLX
UEePoZAt7Fc9Xco0CZqwOnlcqEJfVTyyDyyDGIR5lp+sTHbupMzgexfQMer1FOS8
S0w3Vb/a4rTa/HE/oRpXkH1zhOBxTi1p7qZm5/ZghLxtn9b9mYuU8j4NO50OMOJQ
f9AFYsMD4OK2WT7BUQXFl+E19VDdqbQZRc4i04z6eJWswKH8nfhQwdZSVtqto9gJ
GA6PborhgPU6/VkC7r4SgV98kBDqBZrmw7Tth6s3C3AUvAOOFr0nAqfbP7KmW1QR
GWtDcegnCm7oNHmvmcZN9fsUQeEKsBaL6KD7QBiNFdf/wbacMB4Uydg3vyaVZKC6
JH7tyjKbLM9kbTBs40jJ01TwPqd+a541AUv0UsgPSBlqiyG40u3WrhrCNc6piEcX
ZxrF0+NgAajIuYn9P74s3p2KV40O95e02mXTCMbyagAyjVzlUCNFuNwL0B1qh7S4
YjDP//TU+wC8JUkexlVJjmwOD/F45EE/ZhZGOPX7knH9OiWsJtXNJeqXS5uaHZv9
L7FHF6pOqvAoclo+AE/zkIu54iPOn0+p0+3yxku0kMQr1hJsKZ/zvRrHIqjIFbDP
HgmxMs0JFXteS9aWSFjpo0X/mk37M+D9iQ8cSWREtuYDZnKbplVM+Xh+YypjfBeS
fY+9teBsM8OS1yxN+4P+1lRWzqpGo4ogHlR9IsOjtkdk/C3bgYmtpFOoI7pXUmtx
HZ2baxfhKi1/5D1KR/YcTqWX4Hrs192Rp53rW60LaSIgA/Y+Qgw0qT6mVrwYRT5G
HFJ/CexU/78Xe+i9t+47M9DQlvqP7muUVZcoRYIEq1DAQKg0u4Ns8TIVwHVxJ819
lZvmppWZ2LR3BMl0/EwsPnmgLbNx08KhDaU2W8MRiOd0X6F8jvcW7V4AGX6VINkJ
IUvtEj5CRtGwyX1A8EzzG7SHCGX1b+AZpjj8tDMdWpE3RefEc0BPknkEQw7EmJhg
0JESAaYOcRFg7vJ/Rd+4iEow03NHsQm3MRZWY0padwSyBpMkJ7Yzb6poOj4ZCgoe
E9kC+Ix4/t7aHfvAtH9DNdtb27C5VNwQlF8WZkc3dffyRAX/4IOReuAcU1ImtuVP
6w3mFtLXvOfgpjUS8mRDGzwvxujMUXAQKFrMInk1ni/xUuARxlsQi2UPOqmPSAf2
W8g/OeeXFZ43jyrP8iErVbt1Pu+MpFzN9BPFoW9eRRRkkTmPUF0CX6qC2tlXcdEI
bK+W6bDS9voKdShATDmKNfed6eH+DdoPtT0X62vv0uYhm17Lm3QFCok0FOwF6L79
DJLOxlzcucdpC0R19uNEFUsx/P768c07MyfBcm4G0UjQYurFEw9g1wKvJuxpju66
vvdS5i8ptOJ+gtn3kn5il3OQ/CpeQcRrVLq53FSeLDTC57etWbZHq9ou9lVizs9n
e/8k58YNcys9o/3rBF9RTRKa0ia/ZuW2k0kstPqw3RTRgd77iIdO0JKw6j7NaxhG
RTR5gV7u26fpDIBoxzXhhb1H5V8RRaCZznZFEs0bCeom3jLo6sjY1AYz/uONbdHF
6HXR8yLEwWegObJaxbKyRVT2W7TYxmSCjHfg8fXE+WlBywSMd49NEjdUuLgUB3Ma
5hqS/1WgtGmUNS9MqcqYSSVKgzhhA7Y+l233IIcX+e/KEQkQj1Hac6chFuKywRr7
r2805QRUXwhcLS5BMby+t/7/DVYsEqJAbLNGZDk9t4aUuEtT79Unyi9tww/vkD1q
8Yb1cFSuEW/IfYos79qYfO/1/E7jZqS49fvWto/K2yMs7yckRHAwHUtUJJIK87Vf
bquTDpnukI66OSY5LeWPqmnHdHVAj3HJLyxJ8Q4pM3/Y/olYdk7afrfW2gT+d6vv
MHb5gflvXJYKuoLniWGXjdgZAmRcOn3bfofR7sBrx/8jX3CtxnuGAQosJhZCjLG9
RA7Qy5nKhdQ/4IWc+J3YmsEZWMGPnZLWZBQmNzLqFkq69eLg+LkzrlBDOOjrOH0T
J039r3C62tkCFJKmW5+aeIcn/sSTsvlp9olT40k27AtmoxlDsdQYGlforHNEbEkd
j79hmcvNDNEaDyPGiYX2gpeCr1ofBy3baQnRI5HxVnNVNKofnqcupBTZoltoRc+/
aAVxpnAkaHxyknoaA6hBwu9XxDcM6TQgY7nVnN/nHzyyOx+cMWQecKy/XKsYKPQT
zAaUXOMc5sX/dbeAl0qWufOON+1lppS0SlmNzTDS4/XAzNr0mhjWiXmWEt48ULMI
UCmSXB7QG9zF4VrEN1uYCH42UGLoXLDYbnA0jbCjslQuz/d46xfBq7jVSISex7q9
Kgla2CmtWsoxxCgbvMLjDJmlV68X4C2/Qsqsd9RQ0oNaZNgoszavmpe2WoB9VMxu
KGPauLRssYvwRoujIW56u4baQF4bPh/fnCJ2YiRwnFVaGnILcLrqQdcl8GbUSb5C
lyaC1i4J1u9iWuc2TIFTMcRX+TotV5fA3eHtud1KoDKuOB463hpuIygMdtnV81zZ
r3P411FwX8/M3JiOdPjyxiHItoXAPlda8namsaV5EMaFtE8taTMDzIIX3Lqrythh
dLo/qrKcsyLi8guKNY023tb1WZ/+LIrmbp+8CP2Ah+00aNVoX23x2znxeBZAsTsh
+eJVYsXr7+0E/y+pZ+wR0nHdFHwMjTjiefpasc6SfPLkFo0cVVNgsqYlxa5yDs0q
qTiLKyUYM2r3XZFY8mqciAzgKcpZa/abw3qBn+4nYTYJEK4wif46nyaBAnYbVjZr
mj1Q3eySzkgNxKtyNmMkN5SLxtje7c36he/V4VWwPYOtOYmql3je0MyyPfCAhtct
TAP/0Aft9JaSjh+ffZfcNJgtf8IqY493McPAAYqeeMGS1VFkZcPtn8XI+rIeEWCc
5yfXVuGOsodWgCJIrwxcHD8akj+uoYXqxT8nOYRkvzxj8pdwHSHzOVQPj4d+1A5Y
oFoM38bp8sny3pw27KBupN/RI/a/MCC+fVurCoVc7T+p/4uK+J4GXlu8GlFd+X3W
HPNynPEIqnC5MHnoX9BuB2lUZCJh116R7KJi9oYPf/JU520uZQ/My+UeoQ5lsxGZ
HzF0bq+0k2IbJ6RJfHctd84o9pT/tf9J4N7oLrWndfOXBBps2pvHBJPI11u/O2bf
JgUjBtOP7tcxA8oJBa0p5zCBbTTjTqZhlowHtX7bMCLN2dhoe26LopYtegIBJQvv
YEMGSwHSVGgPPgyV4pfVr68GALxT2K4qKqlNWqsTLUiTyEaCccVWUKkl+jD4NPws
hWRPMpx/tGWUNm7G9VdX3wnBNImWaQ6iH2mL3ZNgsqBrkHjG8zxJWc3YZNlAf9z1
I+xSUZKInfC7kgesHpCZorZoGoERCz+5IHrG9OsN9G5kqlm4X0fXidxHlT4qCAXL
XrUo9OTxNS762yXiQ0kgEo48Ips2pTQOJ9nxB+j9bVM220W89HcMvsEH37aAaIUP
7yYjO1VXmsaMpXwd7qQhE6ESTqwchB2shr4MUb0BzkOMCEqoTZ6Yw/XchnN0aKGd
lx7dbZQlgQRpSB2nSq/9tEaBumM1L4dLzGz4cCSi3vMUN5TJXqVPmkAGoF6PQRsv
5VwTLOv/g95seckVH7ithfbMW9xpJ8jC7LKqdSGsBOtpdLorPYQazUjS7eileUL+
YC9a0q5tBDggcXL7j4+FCUmClzXEEaC74XJhp56hCZNcFfdC8GLMz4rKM4d/AcD5
NDDbXQrZLCP/24P33pwKdvGV0msjiayZbwOHwTtoOetEB86fAXOYyYhYntqCB0ZK
GeuQQ844UWwgvj5nmrgOGxIPY5wQp8SEswAoe/zMUh3bzGBQfgvu1eU5wjj9+x7p
ZuVJWZODD/bLjAwuG0m1T0E1NDKQvBzcoMHt0R0HcXxXXqh4RFyvaHY2TKkL0YNI
l5ER3mOiOYpUPaS1MkfKOvOdrk5bRami5bAPFtoqPv/xdPnk6i3r8Ngibh/0YLdv
QXF9lxOtjLcy0cI/4Sml8HWBf102uNfUlUneaR5fzKMes0gsrPFIZXEvhwaGthFD
76z2f/o+OQZCzJ71OFVQTnJCvn0kVT5f5HTqXD495RDgovQoPyLXfWpYrmRzP6VS
AZMsLgIgmuaHecN0+viWn/K3Zh/jPF0XwtaBH7JR598wlK5qo6O74YfuOEPEkA4A
uc7LxrWtzMEQDaMXoBtIERnHJ2I5dGwXRJ+Ocfegnz8jlNF894jrAXc5Jwey+9zy
MUfjkD5QGUwQsK/gtQebb0YGYMwwr+xYo8ukRzblZ40o2xf+YVt9Ar00Aka6SSCx
q7PL+LwcE6bPXPJ3hd+/EZzPR9wBcIpuiFKB02oB+oGWebzPUEdJrxdpTXkcffGC
4U90FtxmF7+geH7CAhd/i52a9CO/KsRG/XjEWzQZJ1scX40NJRhgpo43oCaHz303
dktuRd1Mb1+ojYXP4UMHe+iGp0YEQltqiWYQ3jeDUqiqU50Vm3jJYvgZRG3Svi07
oFqBo5k0l7w/zt7evMqOih4NFPpD7elerlJlUjw62YEDXftfyDByHmGJXsTZJ54S
ge5d+yms34M/KX1BEYVEbbM3B3ajQ0lPaO6vxjcw8vKq3Vj3CnnC15kIYHSs1doA
MqvFx+WQ9prXBna7lkp27bGnkdotFD1JVnTsa9FDzxlm/31xjpAYc+yZzU+KLaij
ftunupkwELAZdMl82PGJ27Vp5QxipIZWRjmQCJMM026fewgCmypdSqWE0MBbmne/
/6RmS27r4I8H9YemNzc6KQYkKiCnjIR8D9XmFEuQOxSBZLwNJRQBenuTzcJYBW2W
Lx7G+FxS42Wk5lDM+mi3zh3VDCGOKIOA+4I7mil30uo3p1GFNU9h+rGxGjJfTNKF
135eeu6emqHD4xKKnJkxz1n3lDkddiwqj2n3enUtfg/Bg+slNm/Wniarob2Ek8Li
x09TTWca2mI5xDz8nNQ59z68eAIP9e4YoQ0Uvrz9rPU419pNezsIzIiqolfHwpCh
D6wZ9qsNNY2ZzhPY5Q+nWdA6leohKCJihEEi8nTFgzc1RkiRdgXm3XnY3X1aU++4
2I3vgUnIzMbYXpV8fqInXxmEAzTEW4MC/NHdNBzkV5XJh71uaVVD4wQANN4jYwf3
BeOfefXHP0/iW45WIyzjQhsXqzhEti9A5ZNf1t/Moo4Tz8Q0dXZHy4ZMYxX2x4CA
11toMk94sRDO8aPrFpKuei/JSOhp0I+oRwJdmzaB9NxgdxGmfacYxr+ePL1Db90c
XFR3i+sg8yigoQzD9FNgrgphZOH0ws0CtSN3tcj4g8VV9IUMGXCVC4DfDqOLcwdx
lEX1nf8C59Cw1Uwbi56R5VKbp1KLm29+N1Dz5f+bUaS9/AKn3TzSPyaz9Vz6uE56
9zzswlZIpWrs+wV8KoO5BTm0rMuDvO4VjEPo8TXs3CgbmFpgXJEmvH7QhdABcbrD
X9BsHU5bFTUSYvzjyNA4WVRdjlFioxoCyk2FlWUNE37TVbp+nAOTWOwcBHezEf00
kor4D5ix555UPMAR7LNcYjpiUWbZorP8b/8EJGqMR7kFlmzAzzSLJFVaVPz1qSGd
Klzepih+2eTCdJUsPqMMMdNqzlwgJoNDJdd3GYHqPzL5q7LAxG+jS42Ay0N0Y8MQ
5iBFqP0VWRIqS/ZKMR9jp8VQC2aFKbm/U0y/MWYlz+XyioxXGRohcuEc0GIAlT0K
/0+z28FCmrpl6Ba9PejjBPP5PTP2kl1JQBVUsINefFDz5YHiqqUoP13Gh7yq+GFq
cLE0fvj5fgIN9kTj0U4rbSLjYI9bL5Npf6i2/p2LUA33OYXm1W2ean1EN6Mp3D+R
ZY9wIf/CaYc+zvDUHXwL3RxxQj/IfpQlvnR/ZjD5DDI+FZ2YdIfOSzI8f485KZo3
iLdKqCA+AKjEGet3+WY+lxfTdY7NT2nyLrW+0T/TncVl/LeYvYi2MjlZj6pUmaYH
y4hG/aYOE7rSEG/rfb0eB2QuOVVA5edIzVvSfmjJb0RYLsUqOhvda22ecahwQMA8
K6uhRkqE2q3JEVRsXWUHQ48c6R0kzjZaUYqcAX9wLG3JoO6BQotUY+19Ol7UoYwr
gT2EVHfk8dt5L/cUBa2SmuExyD+qHM4h5MmrH61qhr3oi/RnMMFWgHzwKextrAIT
+I/8IQf0AfcbiASO0CR1AUmz7RRimuZNYt7SlY8D+GKGY29cH+TTZOci2C2HLxVR
KrjP5GDJACgRLnjFNCqVXH5qP2zzhzP1QYKL0bIn56gFv/AfQEEAG2ebzAfdY8m/
Uz9xCOxbSi4XPBCu1xu/Otcm+2uII7zw9pK9M+K3OIF/v2vbzH4bTd7aj7XCR95M
Su6vV8rzgDkwzG/01+URFFeRzuWQ4eEMyKSJ2NE7JT2ECKe0r+jKeKO1ty9KimD+
1Tze8HQcjbrNJtOsvsEnYMN399/7uaGI9rkJfHUdDw9a3XbfXmJBzYCmlDpaP1dF
GndbmUvQsbD2umonxSMwAmYXrRyH4LKP1rnaDMPEPMMl+I39gChLshXqrIVGNlLt
oyo4AjGf0zLsxs4iJT5xjH/La8+7Je6mrk13/RltRD0D8c+co7T037lu3GrPXICe
TdFOVJzdGkmgL176VlsuN7dyOcYMLT58H29N6g4bWFraYA5RgVnvP8OT1fRhbvud
6BCvc0Xc6/itEfLNW2rAd9bFpvnHUq2RCz3vJyXt4Q8MKX7Q1NGyYk0Vsk+KaYRZ
Ak6Wt4uXC1GK7cIk0jHfJ4sHSyf96a2f6s2AZNqcy7H5Wi2ky0iGt9RT+idTNIM1
z/LPgdXZ0g74YYouNHfRc9HAjEQeOH2m/XmKNAL8nvsEBGC3SMqJYMTnNsON283G
DoEJicuJhpe685JlEz1fiFyk6982PdZt+bL/hVnHJr3OmOo4PvGRJJFe+KEfNBJw
8Aws1jwU5e+jnun84PLt3WBSkJKxE0LppdXOqmYaceEaxBTAc1yD/ae4lA3H1Q3e
wT1ddIPb9basCoSAIMUfU1Qd/J3hiI/nv1viIV5Lwvfgg8g/RG9OgTtowo0dqObe
vKP9/GPEgkAqMf4fuRYjdPPIXRhSxAO5MoxF3KW5w0ooOE6jSTVGf3UCSo6Er57w
PGyM81vQworkbsK8N58yiXP9A6jlSO3NgIsNmivJPeKXN6i5vKRD9r/RxKcbn9ec
9kvhJLIFMA+aK0P0d6F2cz25Ht6nsr6cD7KJaN0AVbKKhKMLamXYWTrGW/+JnsPp
tuHYZ3/lgkNUrCTXP9PP6wlzyY0EbfZ4eoXUoFtbG0BOaZ1PGZvD8pFjO7DEi0cM
5gLyPyzhw2RzA7G2TJXeH8DENx+IvSgCzAOVPw2PG285mGlakGZTU+N8gyuVJxRY
P7ABTXl21nnt0IuUwExk9JrbdvUOXe3CMl2+W501fvpjQaoNyQhqvu1PqiZmA0F5
Qdappbk+7FRaJUyRkxJlniGn5UMu6Vdc8jUOJnR4gtl4vP6UfVzPNEoUV9C2Mekz
Ghc+Hrj12jJLjSOgKQc9ECapIcrcG9PzTjdUCNKDwX8XKaAh7xeXwUsHJ9bAkIRk
vZjNhPyQMy+Au1tW+pId4qVXh/1NQGCe53ucCUEN1XY+Ti8EJSfgE+B2+jfOdBhp
y7+aBBaWc0u3P6IyBJ0tpLTSuOuSVON6B2E3hbC4SuS+BwY294e2u9WJVeOTbsoT
TCCNBbB94+Pc/CspO60j3H4igOR9v9ZSuRTaMZZ0gOO28YgEweM+lNy0rai+8zEi
cr+My29LI9gP1BJUlV6IPjKJ+Uk6ETyVgidhOGJGUawvbCmwbi5kDu55FdPYID6i
Op/csYQ+s31ls/mIxXNXijobqKAwHv0YD25zcqBJ0zCeztA1Qnp7DVf9svniKlrU
NBOZ5nks+8X+QVFHlOjIy1qjHhV09Tp+FtK6iNuEDCDULdMM4RRxIgoHhil0Cfhq
AVEqVAobrm/4lZXEMEcgbuz+i1FtVHy77/0qJK1xdD5KRKJoMsXz9JEfFbowwJ39
laMmoxJijTIQwbleLeCtMz4ZCFoDun5ef5fKkC0ye1aKdDA87cJzpJQbIty4RZQv
3Z34zWuwYYuO/BxYULqEqcsbBYIqeyR5o4esMJql4EJV/hoLXVkQIQnnQY2M5w0B
fMcFm9ZI6heMA/yZM6A+MG+k3G1ADe9YAcWEnTDmrxSd+IGYvIqEuEx93eZbxWPY
5Ga1sqpJoe6oI+u4tvNdw/RpAUmcVQeXAiUk5qTLhhPaOmW5uiusOq76ilMX9CQ+
me6f+g8e4rqS9zH6VaHaCz0yd07ygOzHkw7zJrQEx3n/SS9FRATIjBeKXv60599Z
P10rdcGJ/wcDAMuadG3/dG/2YqCQ0R4VzvLE4gKT4JClzAyiiLcRrnCWg9h9LtNs
YSb29xtrmjGLfNk7i1sQ3U3RM4sTR8M5V6uJ9lKmMEne5k9vR2ADNeEG/lNb7sAi
B4aMlOmJQnQ3bNx3377M1SMei+1fOUBBPW1KZPVdHoIWqWENN8x2u3cG/7kPQD4b
dUaNg1S2NmRwnoifAe6rUuvur1fZp2e7utiM1U3hOtB89msjSRg5aFmG5L0ObddW
+zcyq/uoqPQjZP1+qrt2c7vWlNnQFeEXlFnOq1NCY6f32yJv+ymzks5H2VYr1kLM
T7acMoIQwrtoBE0tG8jBNIekYFJEAsV1JROrEo1Iu218pH69W85k4zkiIp6ZHCHI
iNrUjR5Z+hOvHSRAOMjEMX6s+j2ZkqQYPBN2cRGG0AP0Gz3rGrKjSKfmOWxwAfOS
OZlv8E/9OPM2DEW8jC9KMJRuXM+p850gN3G3INGDzPRK94v6Ak0xmTxSw1f8cmZy
BbOkS9t7sQcSOwN4A3DeKVMfc741yJ7stDBvZZIRHx5kLQnjt79h8maRzTQkp1g8
Y+Poui59mAE2ZNRahumcPPDdzgMEKAawxWnursTwOsoF9TuwTkhVETiAAoFqR4a+
skpCslJaihcYZmrJoy+H0IScvSFeFQMxYAUiOT4V7DALYUp+CK78Yqp6sExywMm4
E0PwWBpwfatzlwRiRDLBdl2qVlP4N8VAGYJxcMHDdUotu3cKo3PVd68Xm0AMWeDQ
NVlW80Lq/qGa3l4f0WzNlAKrPYeCwp5D094WvLV++2U8G6clcc3PbuhSHrCgTXBq
M5knD8SeYoQ66jHkAyUtFfX+CMa6VY5JgAgjEDVepJ2ywXOlyYYv/jKNsQMjsvkX
90OMvckko2iaSRR011DDK5gHR4qs7AtDh4GNY0pHIx7hBKc/5LZJz6vt2E1EyXAG
Hqs7XIqtSwK2GuZ6s21wsoj8d5UIQPFUBZaJQ3WbyYyC11JXIb1AYGpxigyoNAjr
fwA/vac83e0uNzqsL+MGuVuOLph1O7I9y3z2sY/ZIZJquRK5SPsAEDytvJSTvw2b
GdkRQw1lgjJXhzSKU5Q/fiuWjxv53ssIxQCYLza8sxvEabM28TDnTFiTV5CnN/yP
0m0pt2pLeaWBHzdBK4UHuZDRRMtn1G6YG+TJT/8fThiat7J2c7+5PhdnAfl61+rl
XdsgfxXRl+M/PLQnOIw832wHzWPS78ThmApe77lKbeSl2FLgptJlutFZRF28uRH0
4z4f/CMGScutbZ6lG4vCC+xMd6BAx88J8LVGnQvkek/wpcqX75b40Ca3O/FM6G6k
uopqjBBNSBa57QG6l60IYXOoNqorhZ+x4hZiHuVWhLA+YtNnVJnozcKsnWsvo9FF
wJsrvGLeIb0lFQtbOUfr/R5B1z6udtjDzwafYBRGLAly9GX7lsS3O8tfUeR3N+/t
mLPHODDH87Vy1IkJhM6VF6Dps1B4bXKfms+IvrP4tYTj/EX7mdUlC5lwnqfstb/G
VbHMT2+LWGpz3EajoVr/J+Ys+0daS+Y5picYbcXuCfu9IoOKy+6EIe13mBbcaVz6
swZnsJo4ZwzoBYlaM0Fm8B3JqftoEd0/uLQpEFDJ4/ggDiLHq5/eOVa6gR13AlIh
w3VdntAY7kIlcy8PzE2qpiP+3kPM53jPJZcTtH8fiAnweXSJyX3cWF9WiAiwv0Ky
8bzizueLahARc/Q41+iEpuW9vBE6TokN+3sPv9r6jjikWWNWSjQdmMBv2rwmSiun
GEuUYvTlvsVfri0CE0tmkdsfJbOkvq76FgJbgVmb8deih9eJwGI0eit1WZRqXDUj
BLBDBjf4/OBorf1QNSEtbHOg77p/mC/L9z6h4HhxzCUAgsoiuqgKt/7A2ozXq+TD
JKD8BwnS9LbBISFvJkpON5wKDkb5zmzIzikzl0GpAsJ+QJBtO4/NJxVdxPd1QQ8+
tdX/jhyF+J+6r/LxtxEjnVisYM3MIy827rM+egjCspgUL4iQXPso/gNxxkG5pH1v
CyfccNCHPkNY2CzkyzjnpXWKqAL3l885ic1fEPVTfjTpmBEZ/jeAKEiL8anrHBM3
e8j4YohPQUtunyNr6JyQ+MWZbOx3KSM8ByP1OUj9ZrHTAYrsE8c0L1BI8K6+Ky9z
EG6sfo2O2uB8OpAIGO7IwqRUiVyVjqfaHrXSHN4EijEtaW/G0Jyj+A+EAIGm0yLZ
A74rOXsj7njEVKDz8RQRxn5y0cBMmtcF5MIEQ3wS8SyhGEHglFZ4ZJAyVqYzrHwg
HUMq8Qq7ptNCV8STmsxbyNNots+C9X9/D3R3nGf0B+L3wLfhEM0BxCH24JCNPcGw
6eRP9qd07vowzkQe6c0CdRrBfE1xVBM8DNUOxvNE4j8Pfkx1+M/WcQrrm6MZPad7
HjuyPXeswR52X1FdYsMnmw06H37o+Mn25NPXYemrmrIED/nFl903vgEmBCTRFlCQ
tGkJ2oCWdoRsVQkz1YAZphmYLvwAOz5UOtplTuujaqlW7S+e/4gvLV/8Im+rvNPm
fD5Ex/FniefrWNvalDB21aqT7BcOGRUWDrWoyWxGkZgHZV9dl1JoNNHntak5+Ro8
bV7/9QywmD+3iotI/s/wqERz+moqWq1PC8Q/hAH+gPuA8FD9GOjitHr+9kTReGrb
I6r/4YuzVDNF5WkNT8r9DRF7FrBDXf8kIcj4UdqggGLmVtmh/g3lIRo9a3xsm1Xx
50MBvtlwiMlk0uZq20UfCG3eA3rYd0CkIev85FGx6zI4W4HyQH1y41M6MHRZ80PA
RToEHilWSA62mSiHJC/XAcdC7c1WNSCjr0dp02dbMOL6J3AmYVwfN63lTPem+yIn
GmVSbe18Kjc7jZdl/BG4y7j4fY4AZtfNezVUQ4bKPDKRx+o4zKAqlWOq3kGXKRGK
ge3ZsXFVGHpoNu3eBUaVaHQ00pumsSaS87mMMpLScazE6QGdQ3jswR6gl2VAALDJ
QoIhj3kuH03dO40rNpJE4TUQaegOYzJ9ZG3i/tUEyiLut5edDo0q8adIo4w1O/rX
dOLeTS/TawSOtZhe0hcfcgHmySVz6ZNu2QbKg/8g3taK+/MRcND3YfuxNPzX9kvD
63VsPozdlYCPpsk2722PLq5V1nRqzaCBJdRYTMXqY11YI+bpQTdS5d4jYzPTiadC
iImSWh3TfuF/QvhWm7WQimHGODyMN1jol/QnbAoVI2qd/+UM9PmLELaiuEdMqCDK
fcIzbUE1QxDGkGGV7DV5jZxg9bwbFoErAPgxwNzB+pyHH4+rVGH0REKSbcx66qhM
Lf0TPazrzm93KKXt5uMjaoVa+l68e5WVzFtPCkb32Ajmbag0NYxFsc5JyYOj3Qno
4EhLg1yqJ0Kpe5KUPk9t1TgwVBTWkrApbf4tr1kN+zIb5LL0dh+NBh74iarg1FU3
rsb7hbHgbFyU2U9BVdQR1pTKg9VcV6NZBtahQ1YnD9u44+efBfNkGYQGAPbiveWZ
/CTwEuWIoghyueGtg1rqInxBvCb1IYoOV1dNzXyhjl3q5LtSYPdr8c3hxKpBtx7t
B89d4lgpM02KBZHjYa7eopMeilmBkPNo3V+jSmk23ad7ZlkwNyDqKcgooF5Nlykz
iH3Pbp/geFtiRI6oIqoBVnN35ixnGyqV/ffmaAZFbn8nhQIZgKqK/jy7hlOIS0E8
W/Kzhme6hlAQsox1zWVbtjRCO3VV6jPbBmXLYrVGuytcxWwjTPfriWwzhRB6AtXh
paIAMP+6lO0NcfocsQKVG2PDKeCQvV6iTFeO2YvHaauYxCpH1XBrli1+Xmn/pa9z
mprBt39uzK1d6VVYxVJqm8tL/BLS1MqydTIoAtc7ORwYWXXM3lKZ6Bnx9TsfS+y/
GVnddR+SA9hRfFsMa8UgVefZwjnz2j2IfmbaeCAgtNGDsp4SEf7XK2lXodd9piuI
RvgBj5b10UtXj1VAaMQXfJ/sbZinopsjHWIkIzoGV/WorfEpk8arPO/gL6gWbcnw
0UAAMxhLnqVW1QztjzGqcTveg7/zyjeCtjCCZYXhQ87ZzZF8HPvu1oObDdKqRvN0
sOar7Nq47xSSyB8Du2CZC09t8U/X3sZrisKc9Z6oGM2Q0VzfUAstYsgRQAjOSct4
Wqb1Cv2N/bTAim7FA7gNy24RsmHUxkC11Xajsww7Mk9u0aIJeFxkK+9DU8ccvAqW
1U3oUsM/zsi1SU7exIvtD3lHZn2C9yNqfYxpX+mvMWAK7SOtQ5YFk0xI+I4Ey/nE
AE1SDMQscihoq2f5JrwSXWnsiIAUl3nwDC3rR3YoA63AoTGTgiFGl1Hn4vyRs/G7
LPO8AOIYPoEN7It2JkLpEjUSaUjFQBz7BZriOja1GuB/xrNzhclbVtfEz2u09ton
cGK3osVF0mzpF2mYldkuNxGOYqtvIfnM1gEdrElTE7YhOUyZkagdq4K1vjsBcDHy
9T89EXMe6eo/4kTo0pp5zXtZ/MbMLe7xH/dSDtkW92DRx7ntLK+6oY+2IKYWIQRd
ibqzJOTpX+/0nKHqfRnJZz7PN4ek6yvmzV73T0NYbUpSh7ufA24bv6vWOKKQTDck
MfTb0o8PoPTC8Xgx2ueNt2GtmGEnkYN203l0E2le5K5FPXLhar2KTqFR6o74WiZj
Yd7G21qa0g6Xv2r2D/ZaR7ldAEimht+2POupeXll1DJxfvRzz2ww1itJ/uYDTeEh
9Ccti/OCjvovZNwHaWe9+8RYKwgJs7OgtqqO3Ah37ERbKH17W1VrISpyCH5briGe
O+zES1gL2OyR6CRYjk244zoGQv7Bv54BVFfT/XWeEYc49STnAlrv/QowYCzikQuz
GODqRgmEqMwFvI+K9gMMgqsj4F3dLh6Q10cVsGdkCsf04la+F3kvfhVX2l8ssdEr
PLCtJ9FnI1266JjfBN5dHhRtV02QhszUmQ2iUPphlNmiaLOZMSUeDeRAhFpDOAo/
EVbUf87x1eJxR5z6n5VZrmrhhCUwCAPVzC9r3l8yR/Z+GM0bQnbOV+BGUea6nEMP
VRD4LsRqJWMkH7zk1CfoJtVKTMGHDLAhdBeh8YkF9/HdSAYlCbFR/LSHTd6ffWxD
ElNv54meLv2UDRFvKevNfmF64QtIeGJ0Y7YmStySUMKfF1KAOFfAtB4PbGnK7Lof
qqK1YhOAlzqS05DpL8ccjSLTEDm2dGIPnknw+aclCexxmcp7BGp1jZ4NmMZ5Ng40
l6IRC0bEmmRa9MgUn0WKqZwd9PzPenz+QPl3kEcIj8j2NUMh/FH34KOoIUE1BX2g
b8fhAKJNSIdDrYIEJgWU654PVBRKunCbHpja5C+Wz29Zv9/ueMdxx9+f0RSD8T9h
AXJcPaVp5It07nbzZ0+TkhvYjuAot5wHYnBpRlxXz/hYkFDMZh6ChlBSEqvqh7uR
+BqtdFz7Uec6FwiP2gx2o82lflyzd8E4lqVJmwQdw4osDRhpeNlDqZ/fO2xbEaRq
mwVKnTm4pNDlOO4XfWYflT4YPdezSOwq9ABY81yUH/uOMtNJVCDdlXYhF6EO5kwV
tMl2x5IoEhZJaGySe+ahTTw7f7Xe2wzlcAG0RVlVOohFvNWuKyY4sKgsgguw33zS
7of8F0KdH3zDbIuOuiHRG54ZdZFFdYNifhcq8gLRvdMYHtV4fDYvJ3jN8iaDUEVz
IUve579eehTJJoy8iAXM7F0VgjfeK0NMOlx/H8F9dqOvBzTBXNDE1Q6ThCQOS+Xs
buWBc5hfhUA5d6K8LJq4X1lCZ8SjkJT/SC7q6oUFh4AQfSc5ksd8PQmnX6GK5MEk
71jR8TZ+8Rnd73hyKYNd3qu8PGs8mSDgonTS7E/6uSFASa8H1rLzYx0S4HO9rCcR
aW9M1Jr9y3b1/zYw+X5k/NBK73BftFQ5mfkbrFcgCW8ECH3nBWPfayWBR2UbNHSm
t6ZOj8GaHQ/p/QuW6/ES/b3tYhLOcScxM1T/qMXbnNohQlobjOjAd8RkTh7cgVSl
XF5w9pNupy1p0KH8r2u3EbOSATxCpQtj9Sc2EqTJxdp7Bvu9eUoEr9SkrMQ0kNuv
DCMHg/EQclSoHAxKkND9QBaboyAuJ24pyCBj4YAhTTU+BhqARGpbIdSeqiBjnNCZ
HmSeKJiAvjlbkSZK+oLwFXRq031u0O1/MXG3uQ5vidZsVZDDyGkd1DJm5pgRz9+7
idrUaBn/7N3e3QCbNsPkwLGr6zhhBemWn3fAdhQzPvliLWM2jPTF0QklWBlLFgsJ
gZm2lY+h0PPeIgPC4/k8f4gmpWz4DWABrWVpF78jzRfPMLH0f4oOQH7Vm/dSvXk5
N0WFhHsibLVEvTshFNpQm/P3Mfge0oKm46tuhBjSGbHgLZBBfWL0HO4fYHLD/OwO
x3W/Da5BLAQAy3osR1Nq1AaFrTnQe/aFWtpHWQFxG0wYzF1SAzOInXDcTK2EQD7S
eaH/yURjeI5FjrvmVdGTI9Sc5Jd+W8L8ak9qhHbjCXYjTWvTkvIs6Xm0oxJsvJpk
J0AIdQsRSd3HZx3G38b71rEsBUsFlMIe/5LS4BI+MMtmXmjBFQr/glnyZGLNobl2
duDKXAeCy37YNc6fXLI6HMYGmkuHA9kkAuwKjLduqXIIBuJuW5hUL07hPx3lZT5u
FtCrvzTLaVFgjG1icw/MXHmPOn55BpHZspdgmtLeULmt+lbRHLrsAw85U/oLm21H
e4P8QIYD/246y9xx6M+9EY7lwKUDVjOCyh+pj0vvsc1Bcg3Pn8ddw0bo+81baloS
lOUHRYpDd+L24xsL3BGxiDFvDOtzDEtgsJBEdXtJIMmEUJ1YDTzfMlSWTNRQZinR
Ny64qdYPdM2P0LhM0Mg+M6HB/qViMbLXycVV8KlCTeFKPhuM6FWM0WV2frX2k3KQ
T3MknEEBtrkuVySR4AT1N8K3e21ttf0QUdG0FqYJM4/0pm34ZcatohfV1eFvQRns
XS3gwE8/VPXneYNzqZu9Bk4c0HYzK9umWlspiNYa8Q0yLwbLeMabUwmDbpreISrd
BSyPZe8PoX+7KlYS93WKTm2LI9yM4SUMF2zyPcaZYYH4JxadD9zCxLE/UWtvJpLe
MZ5oGD7td3+UYgseQv6N3MjYUoU7/fdy6jyx02mmIM+Me7l2+Kmidik1J0JmGCNm
SzRXFn3Tc9CoC0xht6IW2n+EikLip4Fc7wA5mKQDBFOyYBbWWuIK/U5sbauNdNqY
5BBoGmULT0mghTuGbCPWMjVVUgkJ/m961N97uGIIm78XRNq09tTWKds598cOJm85
kQA0DB9UqaXLhIL2JWa4HkW1sPbfD09mhtR5ybKSxStO5CdLu17NpMgrUcswWZOQ
D/ougmf/VLwxymbiDigKc59fC765nywBjQ3zP9hqtRowpfWx6ab5zJS8LoImkM/w
0SeasDfFstGFRDQ41pNyZCActLwDedVF53u2x76VofMIPzN5IsBl5oO+71ibPTqf
NsxvelA/huBHwevvIpW/pfhv5QpXoGZrYfsLQBy9lQVyWVDjJzUFa6CdgF0WJQ6Z
Ws8yb6g1U+M7ILvK29+c/kjkUPnbQIsGfskAk7Zhau3IrvGPB5UEOpnLMunwo4VX
099sOtj3uTikE0iRRULQaprVfv49364K9ZDPywQMh27JaH6ZVyfb/0prqvUgAN0x
aKhGQnOO9pn+nAlBW29HeComw6Uh4TkOiz/u+tpgkKbPNnaTPy2Bh9jCfpgx5zry
jMmTq6kyElJ9zPAkEg6ubqPGtOzVKPSDAiBVHlsiFUTWul1MDrSJlmsENX60A5v8
6ciJqyA9Yjrh/+H0ef2T69ktrh1ofO/rTL2GPJWvpnT7jH1vJ4wS9e5wxfQIW8l4
JrVl6TaXLDOCCGxG9se5C5XD74xBJ5TAm7K6jvyMj6MsqO4ISCFr4mzzsdVp7Tdw
vMsfRDD1hXeTPyhTQp1gNjxujoJpN0kZZ+603PkmoVR8I7EmA0tV7A2qyCze+4kE
DasboNJQaSBtTNDGs3DViwDsKIpCbX7kVUYY08yJwUZaFM930Ct45gubAYBPRQBG
fKsDJX5hLzh/PNjtd9qKPsEYwvBn1p9VdDzSjD+RpvZdXYzbtZ/vqT8OBtpM+3EZ
eVT+lkQLo0MudUhPf8n1Vnrs2dy6PmHZjEdAieGv+dEpwq6qkviPleAnKhOE8olp
5li27LR9C8nlmld+pFH+bMVUGAC04LcebjCSPTjv6Ox6VlPkb0kAS04uvpwCg7j1
bdggHkzzTMB8uJ2yX5HpUm0Qrwd4sFxzOnWgcGPJT7dLEPflfn012pAOUN1u9bPB
EPEyF+EWxUvaFJ6tnz8go16bWc1CK+3X5tmXRjpC2IQKVHG1Y47QXBCTY7+uMvp6
uLZ56IS3X8sumUEHoqiXN5hyAwutQ2ox28FRBvnAvNUyIX9OC5NtVr3i3KtTqtB/
saI80IJSL/IbUZSI/q9IrJv03PGVHlu8Zu7l+DDNsjl6dwuhGOjUvLUJOvIIkx2t
cpCpeAgbQ215AsZeD3Df9xNOaXd0JnYUeRfcoIgNczEgNX8HtSVeBIuQBp7M96UA
y9SvVrxWu6JGKokWpLwkWxGds+T+RpPybdxyym+B6kw+6+XgtA/gJiM8r5zlHGLY
7kSCX8OrAphX6wMxA76YsIYBqNENgARV0gqOjHMVM4r2OFoC/HFjS4QtYlehxABb
pef/9qRwJMYRlKwBKZMEjrfoC07d2rMdYgni/Qv8rl6nn5WNCyiOKKrdn4qVG/7l
dju/0CdOgi/voBx7qDEuDCvEaow4H4fpz51ad/OjRKmm6xTWdWsswve6DdgX8MwG
ey7nn5ErHB9BCfbtDKoPjUhtnd+NJUe9rVhNzigF4Doz/hEC42QXsSp97/8RrSYL
WTGXDCE+/8niy6fdEEXim9P84oVSxA/GTJGvNV4MdSpWf6HHT6vr1SF7t7LeYVeX
tFjOcrbilEyIn8q9r0E8UBdRG3lYUX9hVWv1doDN67oXGU2C/jrRBZHQoWETZ/EM
2H+NKgD3m6KBC4biiS5oVWdFSOYfVMGNELnNuWhJRFuxZxDPempT6nr4GX2FpIhz
ufPVNJ4+YArwSDxYi+1gDKQr2yYKWYKYEy6J35p1d7ZH7pWYb+4mdfvGmTnwHGe/
F3UC2LSEaoKLq5ayA2s3VDB58BY5DXfmQRonwFPg82I2bNXwIew8vw987lTlv4HV
ATc6SCZtMMH54XldLH3pg/kWQiz23hWfSesWwMEmGN5JSgQTNo4RPgo3eA5L+FMQ
UBVdJIbAKWrdVOC/ocrJ/aR28OGc8Sk151+c5ekzb4Siuvcfkf6lvxMrdFVu9xeo
WhBVtODHTNQk+2+T2oAJ6f/8rcxoGHCv2FhKiYBvZBuEEvgPJ5hGv/NHYAbDpIBM
a8Jr1FxM5GMjkG++o6xio8TIqJLMZUAJl86p4nxz+77RjAEiquNTDhBPjwuvtayN
q9Rg/oUOXc3b3sMUmLFgOnxPSIR2+DkLdGasxCl90zo3t6OoYazU62Xj3BSE6/Ua
5kinzKPE8ZztckKbn2AS7k/xdAjr13VwsLiLANJhHXNkfF6MaFywWU/uXmXcgjiO
sF2AhEBfJgLVCMMYpypxIzJSuWuCaIwkxdOeNXR8gXcjmLyRZhpIpi97YcWXfZ/6
CTwpX+ijM0uRC59kI4mYiOpkuYVOHWKXgpCXs6RFxeeEHK5vYIzk/e1J/DnS5BZC
RYQr7pz5Fit5ivKrsDm2a3bu4V8IVGObWLFmaAAgAeUJKDmEyeCwv+4Sygj+XqpB
dsRhiucY8yF9cVKMM9H94nsHqC1heuE7WME8xmEdvGxoZFGF/sLPUe6d7wtrKfa1
LznYAmcS91zYDEj5PQ7g96JTk6czP2QFKWXf+yRvLRYfuGAn7bY0CCDwBSCLgEZX
gSDWfbr2ryuTwByeKYergLM2wu7K1xnGKs4ngdU7yumgy/xMB1CD6pTagUHrUHM4
ZkFSQ5OK5s8TdQm7EYx1eK595TXC/TgHag6IW0xJblcivEDwhV3Hf1clGb+LNRft
kIxkdovhl8FZxuR+6TQTF+xLAOvKYeRLC5/444GMBcvn+3RWf6UPnN7GelGztJ5M
Vx2ajg4nIz50lUOAhenOM5svQyswUj3V1Vup4X3sYgIhcHhhBzYU+PJO4gWpl2AJ
TTPD34sTL0LVZ/7YRetgj+tePiCo7COu75mQrJPi2P6aKcp2Aa8mU8Knh41NC32O
F2cNW9qoiR5m1wxktJbIJbZ/BBLlCjx7cYWGDVaSJwE0W9vUXc8NtmeUeaEYpBkI
cyA2/yczZhOydbnWD56tRo9F3HIWzIz6aJivt3FXrvN/QV7PwgPxnIjjtIkSbZ4w
4doSlME/4iHQIoVV0Iatkec2nATZhUUafie2AKv5NOch0uuWvxIsEIZfxlcnQoEo
Lpm0isahJSOj00p7WgEL92GhPTJUmQ1nvSQF1CFtPDmXMpPRfzDidkMu1ydJN+yF
namKtToVdNsVNS+6mLTi6Wdvev665R5TGEctCTsT9KRIkRLtbYVKUO9TVQ5bvXnU
TNlAeXrQNwgTOsXklbLjRfkfIZdj1J7AiMl5lDbO7J/Li8+oxz1ejwrBq1DNPCDc
hszH0/YjmwKFunC/pIX9GNFdw6H6oYtYsa/5+wg3QGeMk7ntrv+DafMWHUuVD50C
pSDj/U3snG0WjhUo6yUtfT7EoQHw9TJlpq0tqrdsvHIU61nypEyp3YvbqlD4n6La
NpaaFEd+CG5DXq47PFspgJln9y/AmIGoOtqnHOfSFW7ExV05F22Ax7ZXQCl8Rllo
Lhfnk8kQsOlBw/DXl0DVO4J4PGIoX1NWBa79OZ0ytM1TibOW5wHQNlYw9NeFxVoy
TAndhh9obhpayVQBdB6FGEQaVPEa7PpfcWRu++B7xlAPhCmPPXWJe4OGmCvU4lQ1
oVHQ1t138J8hfbbvYwpORaYf98xAxnsoUQQNbvzmjd98ijFryJP3d0JirUn/+wSM
wocpNoFQVJV5my/ck4TvgubV+GsL2Utl6bhsy8AC0hq6N7LGJQmW7/BoGGdmJ1z1
gAumrOPAi/xxfskggAESDJcYfq4J/O91nGkVGiwbymRefdicCeS3/0njQrwsEezZ
W0vyHL1ATCaSUwpXu58Cj+/s6JspDbXe24M7KS0G6daP+6k7I1CqAgcn7ExFsKwQ
HOlJB9gsGhsZ1lyF82h0aVdCEPzhqKrGnHsNpqV6C330u97W1gaDZBEGfmNDRwcK
Pk+/X32/tb4grNA4lWal5gMEPhaQV0YUQZmz1Qp4iGkcCYnXn7yTeB1Zex0eDaYx
vnDlCW2TyusJFzdtBzPx1lAf6FwFQqiOAMmkJ30sy2wN64hX86i7mRQnFHwSs2tc
ft2gv0096VzyUVSLGTknOJFqMaPN5n+3GK/Vxbqu6bm/aLrFbI94M2VMkjaRKObb
1miAnIefYmUtJ1WU46FG/0vwJbIPowu5NoUdnWmqvWd7t9sVntcWlk4nAesnc5WB
xjWtg08q01lBfl4bt+dkgpM2QVGssPsIr3mLdGcZZaYbl2mAyZegB3yjelypkyUg
cgPe7Orjjb5CfbAY41KkpUnlaHywZoExYN9esmtOxKY+h/iyZKrKGtW42qweNhQm
L9sZRI3pxPLyTWbfrn0cD+5y9cuyRRJtFu7vBypsrDQCwxSs2G0y97gFPgUcd+0p
YHBvVgOHVKOOPjX7O+TKoEOZdeV9OEOmPpa5NF6o9nmN/z00pnIZgAPYyLOaA7BD
gWrw5Wgmxx8tZihveQwTGoGSU/XTxpZ4CcEd4LZpnX+J5HjzPQUEKZU9Nm2qWbEP
XO6R3J8z2aJJn/xTUW4hdQitbAYSdMkvvQ2rCdnw00tm0T242TwvVHfN95JzXEAN
7LYXxJm2nWOjSW38NPKQ+18jrxo3m/idgAE6nnEO7Q0SCRE7EN+G973Vkr00RhrH
ruy5eO7HWi6Gqm3Y9Ijt7Ymw+YATIUZlNyNsfOLp1w33nc/om6McVFX44WJTVOe/
1FBrT9UcIaqyuVt3Odn/ENUiITkGAFm6gc3TQgfTzfpIoRI19+adN/txmzOlPphD
3f09VuIX3CCD5Mo+WvwHPCBcoPLZd0SWjNwUTM99t/HH+eh0cX1PVrm1/TSgpXc7
69AK6yvEGcTZAn5nMNz7hJ5OytPzRzRNriA7a/hjonqX58efi66RTVHCYyV3KGPU
V4ybMxustC89xkO5+cpfOv2Jinbzi5woyPJgRRy9ShBfZN/jLWYT6Isfg4feFXKo
7rMPz/v4P9gGoaV/xLNkfkkPm846Uho/7MfP5wqyxhN/1JibBZhtw1wCaDnaGGwh
sqYT1/IeuX48qQ/APiuEbOA9/Cf4R07+c4JqE7vEsT3du+OMZfEShEXsThifwGR0
0ab5zusZctpWeQZRKY0SMK1pBCYA2RynXes/X/2BepbJYK+qdq/J6TOBBGQr6e7N
HtzFpsbHbPl28mLX7Wydm/LQ6b3DoCuxeBtFmbGqL7EeogCrNf8MId6REnEWO46P
8jmnHOIh5vtViVK74YFp1L3uiRao7OmdAriSFTzh4GGm93vt+y3t6Kh4gO+nKOk3
2MvbgjToM3cjyy4UOOXGjeAjZM8tl3OyXhUpIF+YlQDVB6lZSXvSQf967mA9y0Gd
fO8zT566Hlfin1ByX5yr7QgZBCQvjssDbhLM+8PXZpd1pdnul0MvyCk//4ta8Ka1
fuPzfWN32cnKqWJf5Icp/q0Nf3J712IkRh+sBgIEATwvAC7POeIA5MFtAJ50XK5Y
hu705xZ3j0Ds/LHSEn2NEsDUs54Llko7HRqxlSR3SBPEki5giaU+GNjiEIq6mave
pvjohgOBc1+Muf0EklrdS1LMZZvSg748nyeEyPVzopixNBWiZlXeuPPnrWpR6Yim
fHbU2da9TIp+ECgAmPs+1pZfg0PDVUEDJa7ocV09VUcu6uBeLtJ1F/uIX9y4HIvo
6IXV+tyFnGIen842UdQqz1l48fCFhQOBVpiGgRkhhTdjMtcKdk1kRDspva3DfFUU
lX3tUVwq+z/w39TuWIxC2UJI0iVYLleqZ2UrTt3FhTScSwwrs9NzkSzBCM6nYT0M
R8KC96wcfBvnLM4IGmZ1AclLG3woVK+ZiCRgpdcLoqUte0EI4JgHxJugen1VWVGw
mO3g0XzQ7EJOc/fMDEqviDXfXsBrgJ3mj3Twzjb1zCIj26aoVyDuG2IrZQUvUxW2
FI51X/fosHN3pSJGgavc75Q7rCO9LZiDHbW3DAERj5ItBa19xG0ZsoIMETEjV9rn
nVtf98N15EGow/KBikQXmTyslJ/nCRqcEl4ARRK5ESc64oeqOURuD0M3qgP8wmeA
1lxjBG/B00Fzi3A3YNtGy+o0IYJTzwrwhCYZ4fjjRgIFAp3BikfIvibY5HasUIUr
CNNi1dqQppeSLxFwxmcewcSVMcplOzdBN4KAg1EY2oCaCTiJ/H4+h9HuebHra8ts
Iz3MDJ58j+1jqfUn21ayJs4QAQLF75wIlY3+5JWbkvRUCEsC//P0NiRHSmhOV4xK
8zFed/xdDQklBRZ7ZqhZheTja8/Cr8TAhBH3AZuB7kCLDn8IqJn4e8w5GQD4d71U
nLPur2eoVpvIbPKXp+KAB5fAw2okjg72E4QL7oDPmBD4G/JFTNAeNao3Uug07pEU
By+7PG4LlneU0LVBsU0mAQaRHnWy1dvMnIHn+XHkezX2PyxGiVlkihZQgz2/VoD6
6F3nVK9y1QKHfha5WdWmNWjNCnjdHXOVg7eHoVLMMTUs7yfjtfahG9uBzgrICvGs
IORIStPCOvj2f4ftQWepfwcWijEf8GHI9ReNx+GX0eJB83SNSbUXDnk7P9Zildmz
zs7U6oXF6O2uPi8CdYdpIMrvcJz6D8tHBXaA56m1zh7/pg1BZ6uaUexfv5sO+ft7
ZCTBSR3ccdmDR07DrwbW2N8FVbGILRAEiu/ST/Kq9T6guzCcC09Npz4Fois2h78t
/PiOkw/ReT8MwmUjC7yJVuWRoDBnENnq+9bWG694SYbIlL7Lshh9jYoNsn1kVOCL
YS1l+tCaFTy7VA+V2BP4TSAmUDmXXzG1ODXqmg2vjze7mouHsxrRcpMERVKen8mW
9k+85GriU6eACEqb+G3+gJOCfcy+GIqUGMf1xGLxjcwdSLBBaEcCarp5ixn3TsT2
phCZIiCbDqmhGzUrEHseNjLd2fFhf3eyr11uJyARo+PC8jWBRvko8Cahs0o2gq8Q
gxOMZJxU232deiII+Jpzdds6tSuyo7hjMybRUoE0gB3NqhlqcMTyjG8roIDYa5pX
BaNk2PlDlcXuofIdbUzfv5leVFV20J1XSyRC2TDcJekUDb4lOS7njzzti8iwd7H0
MzqfVQRNBQUt4m9r+PV+6wMKQrUXtrZLdeYruK5LYaQZBZoKkwvoovpRUjGYoXd1
uVeZQbXzctwUxUGUcwapGsqaRdFokzuI6ZB2MEdHb4nAZ0293KEixljn/HZS/mH+
5SAVEUGrDnXLo9iyiy5/7SxSrcrf4U11vS1m+dwP5q+GCFSmDDKq7F3qU6EJox+I
duDeUXSAHGiCbGbJizDwn+21pzNgqOChdWzrnXAEsjDYvBj1H1WtVuh4tf05cd+d
tJtyP5AncepQEz1U8ukaiZ0rCJVz6D+c+tGY6MWVpJMxQvxV/wt84IkB4h/U+EK2
5zdm/lWjMQyYPef1Rg+u/MEyaCMVCnhXgyZGeIG92xXB0nCxvEQrmj7lNskiW0K5
nBc80/zIWZgKdiZInVoqC5YWYqm1v19EWSKMofA6mrKu45vX+NBp0pncpwZiTi/g
cjZWiiR4iS0+zPq9SVARKpgvHelfb/IrFi2tOo4nlUeSN9wEkMuF96YTeS9Iscun
WKHqMzoipgZoV/A9KV5o9gKRkpBmq78t1kJsyIiJKTZoxT/SKMWoz+EumnyrUq+p
sUsN051aza4GV8rGrHGZxawWq7t9vX9LzMILjdhnHj5dMrBJkzyqV9GDvEmN2Xwl
hLXvn/Y371Tlm9/7THpeBecvaLKdgEQijS2+cyADKxneZr4pn813rNJYQrcNNcJZ
lBLZJ3DHaZmdob/WieW94kqV+ELbnEMeFWdHiE7A+8AgemDzMDdCnbyZpITa7P5U
jkano8WZIC7qKttC3eLPGm+8DH1uVZLW2WKXeu5O3qJ9w4XX6AGjtEOGHdVulDy8
GaHQ0kqL3tRsBCYuYv+BoIN+5KweInfqAW0uW5s60BDuwPDAhbE9fegU4bHq1qmf
oI363Ti5v2XhL3Mf3+akd4xMzzt3KmOa3YVRkGkqt8siPq940tJOGQTfY6NPSxnv
Q46ne4k//51MKe4nQuRINAC6Jm/45x16/UrbM1AvXp37JQoNrlfnxoPAe4sKafrA
OoqvXQwN3xRvb7I3587aY1kqo45+OXYOMF39HSvlEPDoScwfo8aNCR+XXnI+i3xK
iJ1+dWRKRcKp7uNoRJ33uKWIYkwENlo/PTFw6EwvB7qZ8OAoc8OyiLJL7KNWf1m5
aRj907MlrZ3XhZi41ps/bzxe25qd0efvymN02LXcNTS/d0uDx7Rd7R+eDqXSKVuV
M+ikhgUMxSusSH9ZqfUcfWCevHVJwAlzAhbKeFz+BspZMlHIu99jf+ZHTpPDn6dC
0X9OPbC3zvPUi936OzXGTXJKmVRf3tj0bZxOpPMT1z7ksMNpC/1J7fQnGJMRimdt
nemde20pltWW1mgkzkGNhY9baoMz1uL9f/bERTz1JCTCmxRT6KbdKC8weCNNxKQ6
0shQWE+TS9kBppWehHcrM9tv4moDqg2nDftFFvnNYbiwCZi62pnETVOb9OsWr2WQ
AoLBUouhVIfV9EvNuxn5Oxurl4FDCa9o0mNfj8RtBwphTtZNuv8obVUQAO/hKViR
KHC81FF0FYVg1jV/Fa3K3mBAFwrytu7R8mFUzoVoRUxIfWF2smqz1QpeFaLPy/XR
cEn2r1vXINWACDxjR6UgSECUfUZ3XWuKgfe6NHBERsU81GBHrz4d6CkylWTHfZLN
0iDR0gfzVjXP1ROA7K2ExH9kRhbJZiZxS10j+WFhTnGEwQxy9mC7gjs3nrpjyZHk
MC00QxQW3NI3tzm7JI3hHk5e2JaJhzXH8NLOyv4FYy6jdvrC0M8YKC4UHTk+tPJ0
kOGDvuQ5klONftGbLFzrGLXtQXQsa7H4KrigHKiX3iiUu1etKyxQF/3Tqi0NYxGR
ubo7eh9BzWO5ZkZFaiHVj1c0nsbKR4Am3x4I1XTJABe4zq4SqhO/eXZz+lRUzZY7
MIpDdm+8PNGs5BaIxObmpOVdOkAqvOoTS30yQwNLJ2nHb1+Ly9VC3w/TmY3TrbK9
cjpdDUV4rhjIuMrlny9VpGy2QBDdiYbT80RRQ2dVO6u8jhjXIwfi6mi2rYc7eeTc
wixKaakeZ/tZiufh/bNWrHufjudpmg7WYKcGJbqnWly8BbbUI4W5hbPQNzYuxzeT
oW88s8xNVs3P22w+moO+6YGeNMwy3efg3ebgqlYI9W6R2sFOeZfgy1dg1p14d+z1
mUjEbZvmxwU7E+2YdmDviEIEUBskQSbxlR7GydpRRJ0H5lhm9xPKl3Q12SoWk1lR
3Ctao9S1rxg+Voru0ssiseo0ykdGD9oFkEgR8RNs4VGqvMNBwptR52jAXSiSprjU
8FhNjMBtUHxeXXPJ4Xy02D787C33rDpqSwpANyUrkwIhAhDtGo4Y2AWRV7p4ix6E
MKoq/eCyxVIvwv57jXsyRdGPjGTsRrJ+WJrFcf1RuZsg1qTR3Qa4sUD40nV+1NPt
zRvDRNITKebPJ96sbM5HP5eTVqVgV+zBvzR024s/Q0Z10rTvdlLNKFqPAvEbtkIl
jzoV4uT7WeqG9OMAJeE00f948wcbVNx8ZnGH0KxpNwn6dc97EQVSVJqv7Xr87PKs
1w42aDqBOCFrEJ8iY5l4JhB4LAWTKWdGqyLqv646IQhTgCBACtCKoj+NvbH4B3iA
s0f8VpVhtC8oBfTFiBD6eZARMrRFLXvwqIbtaFPmqUKOFKuH1kf2zYCTnhbXA+xw
xOodbLQ8JYwGscTTyusloNqVeUkbkbMoGol2G3Ranq51/YnX+90MetOKLJpmIuqD
K4NGhBB4fp4Fz/KCDUJdwyYEk3hXMv9BCRR2u7eKnJd1xPyFcIq9yenvVX/crZ65
rimrhJfMD+OtYTTi9py3H6WgRvV/akoAvb9byiZJ/Ap0Wm2azKnI9nSs6562unp4
dnSJdy3qvviruV+K48mpGH3vWFqn/rIr7SbZB+jHqVDYObR9Co6wBLoZvSRPH3RV
0P39EUHdwP4/MT+IqCn0glx8JD9TOlr2eQqwldCV+XhcFZZW7akdJlNGKCKTEtj7
AINT1Et/6icuiEWdVr8yTtysaUuZMACv0g82Vy47HHdogGpRVLtW7NJTUhSYA+0R
4LJh+s2znPhXu/hNfI2Ne8L9RCU1RfEAsojCfwl8M3blfH5IS64hGuFcXeGrcW/h
LiEv9J1y332SVMa5nHaHRq1vSwtlPpoHBn5k99A+yGROf/8f9FmsubofddC6Yavt
CC1IKoUxnZNjcQLJsqU3aHWgH3g+wIZr8p/WLiGTIOmEhwQm+NdEPZXfzaBbsdYX
X3yrcPZsjlfNWdTPxvxFaztMauo2I3AJZlrj5y3Sibjgq+ElqwvQHYqwbhCa9t/Z
nk+pV5Y3jkneYaZ7JUMFJxGR72AD9DxaijZ5uVDVQ8ya5/nlHA3z9gjq+EHPqMVO
guKHCS231Ma/tLtJPpeU0kMI/mV2Wo3NNigroIGj9bEdkMOAFYpR/APltMMh05pg
XqIoKyLYa/sZUUwT56GZVDLDUm3WoVg8LGi8gpocHkNpeWKNQYVO6rH7sluD33Vc
u07g/KKv52bv1/EeN8aVFxvpaWhcaegHhzndt8CmvK73fb1BnpYkeSGXL9qPR6R5
MlD8Z6WCpctfolIsppg6xQR3Oo588esaJCknGS0Q3tbd4hW4ZO44XpIZ3isgLGcS
nNrh0kOgXokfPB8h3lHFMw2ichX+jUXXOQAcmZ+JmObz2H9qs0Mm3XSp9pKpfnEp
7NqBkJ5NBuXDycXOndzEdta6zg/6fGYThxShTB9lAfTzrYJskttz0y3ZAIf9d0us
eTOx1kpfEEk9Z2RMU1P+zT47R/n9lDJocqRghCOc9mLS4fameT/dqGMhCKD8TfvY
MED69BtObVR/wtnocOrAYsiO3y07SybnwSHX8v+WMQJpiQDIBcpeNV7cw54/duJj
sCvOHoJ6k/LbCfhu1Cl+wqOz1blEuYx8Faq4AbKDrW+Cq/d2/zXxW/KEfrKuGldv
qhypeE50lV2vV6h9MkF8SEweX0N6jlPHIAlPVnIbsAzP24/i8o4X1sjAw225Zqd7
idHl7oboInx1hrnTzx8aKKNJnM+P04SnbbFTTA48RLaQI6R1uHHyZcLkw/eAKL6k
G8iJXCVWLZ7jKT+FtX/4HeDqy5N0F+Zi1JGsWkFOWrOo4/sy9aqum/sKof7Ld0CL
qoAMy9E5ySEE58RENmeSVPr0864a1oNzPQJDODvpx4uzTwxxNpNHL2L0QD4fdkO1
ZeVDPYZKjv4CgK8Nb1H+fQ9ut3eSs18AkJF/mgUE44uKKrtYD5tEZ46w7hpGkUp+
goor4yn94Dnk3kq2ePvRsDvTmh31Ib7tnLJZfkVdUJkBUttGuXcvLDNx3BDy78Oo
5mPz+//5kpBPLcoW1g9xCc4MJDugeeEEwnb80xzkVMGjOdwUJ/Gy5c1e5ALwjQz0
EVV03iJXQ7QV9L4fyvQYAlKg6vAZh59zxKsvO0RZTAf4v8+OfByLMmhOr27yYVY0
Upl+A3vo+DCQFJjDGwbNqBDI/B8vDlz8iLW6OHVq4PR8CV+oa8u+B7vfz1b9rt0w
V4UzF0hbRMY6IfabJmor+NVHCvj30viB7CuxgDoSJ6mpmHI/omI0zj2CONve974x
EELMHREzgUtWyy1PDJcjiUUkKDOAcb8XKdCK8rAhrYCyym0ANIHYgN+s45FOg9OM
BbgMXz3ZQXgX2BmiuHzpTDe0sKWKIxRquBjVCfJHBNg4sEm7cAgVjQBE8SyHnGoF
1mNZvAoQL85IFyA9kDYCuR1pOk4f7KcVNAh6kBF5FahkG4dNMUFSvJaKkihNJEkr
V582qel4XKgtbZwSPr2EtleI3f8MOdQdvoSBGbe0yk0jeaEnywi6jZWYPxl2+4oC
E/BIWUeI/VOLrQnNR04FkJEHZDpM9uU9A9MYsxiCOb8ORERKzQGWL/MBywjxU9qs
ZUoDyUep3NXGSyzX82u37TRzQcv+JmoVBml0X3wbP9pBc/95mWmpLocu/detVJ/7
pZh7bcfOikKnS6NhF6wRsAFcvfWmXZ6HJ1HfT2CbklhVglj09I1MDxm7sx6F8EE3
qEYH0gZzjZyvagr5tBK2Dv5Yq/BiAmgsa0mWR1fYKxgEp8fzzlhMQ7SwPmCzszLi
TRstmA12nvcsrazUDhJ65ofQXotv29ICyG/elICMQFCAF45+KVTez/aHNZpTFef+
djfm0GEV4YKZSkgUGsTTYZMMbel+6EWzAs2Li0486lkMcIAv5AR7vrgOAk5Oh9vy
4qfqQDOge2W265qfN4lrLdjqyILAnfeVgF75+XEfYTq0NJeCnlkMfUDhPWdV8ItL
rMhMB6QSINF1WhjOx4R/QVCAFSOuUzR3x0PXr47jOj8BOdnFbeEuw4TliwD74B95
Dc+kVbW9aZwD+AuFGZ0vBWzs0hMRuZ3GiEvviH1UTW1phSUD6j0sdipaY3InxtGD
PlLCEtXo3AZRMKQHPkivpqx3pbMkhA5zTY+r4KKJNlc0ANvA72D2OtCeehA9/aPT
Z8kEtfxyIexGB3hHPU2O9dsKKUm6jSYWCkWSULx/Nu1CvnV35NLOB6bsZE/etw1h
W5f47xcnQ25QsQdjvjhf3TKn75pEb66MePbxHrvkR8LAOYs/2uZv2Fjr/KQBqNY+
LruxI0CT6z7apkLvZwtg2Dw7XW/Lz671Wmv7OzYzJyeojrjgZeCkHzF/T+Q7IJDU
9IatrmOIUk8mWI2cCKqJkqg4Qgn5P4wPmnvLfGPhog4hhTpL7cHaMWcUENVb9vxs
8LN2kDG7kT7y4k6QayiYlHibD6gNMg9Ljug73y/1D5M5dVzOkQ8h2xnr9yCucyu5
mTT6zmQ6KjyXRC+fQ9RWP8xhvmvWmxkdIM+/Gy1FNEjtQYV0Td9WJh03gwxu/1s8
TVRxrnfxYTdBfmxZAMUKIHOjwVOWwISaNScMqQEb4vspGdz2j4x5RtApg5MVuuh5
v4Xby+GaT8jPMB7aT77MYIiEhDlMd8ipilygKt1WAliIlgc3+KvJApEk+hy0t6GH
GpJ/XreBgw+2oYx+g1IWMD9ydWVk7dW7BzN7skL34lBTHp7/EnYQSF9y/jxy5B4/
yJzct9LLFf0p/VXa8Y6b6s/s05JKIu8YJAuHCfSl6uvHkKUhFd2dflU18MYO9mrt
9AwvZARd7E6OJ6Yv/06qO8BV9BPBZ6VF7NhUdMqpSiAY65n3sZ6yZHe67hqoba1V
ESeDMvFHNsoGfiUtdBhGyiQt0XU/rKUQpzniwu51u4HtSqCwKEXvgZ3wOe6VWzUH
RhNrfjC/cGDU5TAvMg8FuvUYb8WYlzo5xj8xvXWm27b1qEBjgy5kSvwS6hdlSAp0
SceQPHw1AYpp619Yqw93XxdNtZI14hRgWSBBLTHsq8TAiZFsyrar614mpziQdN9b
f6takfHM6NvGurfJgPFYgQMyCRah4holtw66TAQ+9PGLvAmo8I7S8tkhm5Py0UJ1
ae4sAuCW6iYuNllPjM/7cyT0Xf5D0B56fJa6eR+g/hK/1NqQDtLN7kaQAnoIKsmo
fprpgbpHu0CNdSnlaLoT4PDMtT/usqdQNN8TlpgJ3mtCCageQumO/5mFA6wCHsBQ
4HhNTsT3hxIimZU/WLGBM9Mz4Q6HbGs089oOqo5RFL9aZWqH14MH/KRFEQeBxYz5
M6dZ7yNz+YBTJd+fs+Vtpf0kFJUPmA6A/vu/QvlLN4umzfhOxfmqjC5l9VNbgbi9
/cJq/g6+2tDxlaWQVNpSFJvnP6xPqzpFOdi5L1UeSkdrVEAj5FIxfbXUjSSbOKwV
m5cPQmhjJnra2B66pRJ7yMklcAh4hbTT3gTjEtPvsX42Q55Pxqg+RIAz9FNhsbqM
t9OC/SVDmw2l+JXMKEAzrAeGf3JuG+L5VGn59xhRYeVGBO+eQqU2gCtcUpTMIsUE
oZ0Hrs7XzG/PW1rO1l3jGXNh42ZON73ecGMsKYJYv9G8F3axjUHr79nWNCnbsEh6
SULJLwike/AYsyqz5sqTVKgK/TMe4nAmTpJjlcXDVGiT3M3FXZkGETUD9SDVABXx
Doao75lNUky5x4FVxg15LMlynSmzvx/xss0XSwnRjjsiPYKMg7oOwf3jYAYSBWnH
3fua4AjJsyKzYummGrgkXlv+1chBx7ALQlXU9oXRQh/UU+Y6vKN3WKK9R05ErO7/
G1sbRt32JHLBU0BxWXF5jf6T+2vR1FUrlWFFUs+oDw1aYuf075YGIodvwDaOMfq+
hOzAVpLla0QVDFTogp8LLVzv4zybh7qn5+LAmdBx82M0xlM/3P4C7FuGTDUUhFdt
Uz6znChI6MEz9I0Kbbt+KtWkvk7rNHGRPZ6AhR+jsjRspyxHuo91v5g2PwzWRgIm
4euIoTUrWmKG4QL0eBieMYeBSbAxj6TSCGB+Ca5EJ2NZ436kOnjDIae2ExYdWyO2
HJkt9nZaZpgm/bunnugVjQVwn8oCyMgTvqts0kRWK4J3KIfPi9MPIJfxQYc4sGDL
SbBwRMjjevnOuhqyI47JA4lS9iScu18Y9N5kXB1/1Jrb/Q40ZYMDEVrFIuEAt5PD
mjhTFuwbN0H+7VdbZH6jcB2DtgXKKyStDR5nNV2dfqSIRg7pd7UivlJM2NQMbH4+
476Gp3M1aTqYYmAwfkOpqbsN8r1RyBC0jg9BB8NNWwWZdfb6OPvd9NqpLS4J9cqE
3Yt4vrCQ5I/VHRUjqbvDVZQkFrV4uJnUi4sS1TjQrIAKX9dcfNzct0hJ+3WPp+Rc
hbYMt4w+cRdU64jdxvYA7jnPxlP3rI/Kyc5qN+LbAGOOzaZrHl74obWOdW3/O0qb
kuh8L+SzQZv2+QUFWSwSLQg+dcssHxpmkIKTQ7+uOGr4+5aPaQTVJxx7KuamEgZj
UBoJCjmP9CMmvI8G85JFkW5e6kV5IxBb+pd2HlY4pVtpdm0ECqeR0SJFxA08o3fX
/DwcNakIEtM04kbPfp6VqDYPm77Oovc8JdsHJj2rkJumw44BImIP7dCMRyCB6IND
4T2lK3UZLX1NTbEVT6CCgfJ1MHOnl8G3itSviVJSq1PqpTdWWEP1yumtucP2TnuY
O+D9Z9ylsE84OJqqTznhMesZUuzl+txH8GFx77Xb3xn59PJ4de9KrSzgJK7SgPOI
MgQJas32A3adfgaXxkGDHULgg8eU1pOf/upjJDIH2ktcC2IoWIwtNzEP76+r7oKd
7fukv6jBu2rLKc7fYpeDDFZzpYk9hSOKDhrn7Aor0RdwIiNlx1ws7YnHHuPTgs40
C/TFGhTnSTbJoNyWYkWBOMEotAiIJ07iwxcp1Km91820cdLtKM4lEH/PyvVIv2P8
FHGgH162K3dGoClWCCt28uCbiD35ABPv9zZJ4CAF6qEZJ0jy6EqDPsLl7ENh2oX/
0P25b9ny1ieOANGmB4kTNwnirAzPKQy8Mf1X7VaFyR39490JDsnHZCTBt9+6heGi
Bgs7xe5whFswdTMWyvCNniIdflKpd2p3oq4tY7Ps8jeiFRkXQtrBJaSfhv8hfeTa
DEVVLHYzWiFCPKy/Df32WOH98BZo4LLLdJ2G52d8NJuEyoV73CIlXgdRJLfDFg/A
THLO0FbYXhn0v93TSB1/aQWAw6iEibx0Yd8sj1Xp85HXF8lSITyPh4pfeDwnt+Xx
tFHNxWhugMf76HcPflDtoX85MbpRdSn9zMgkjgXvEbNfyqeYenrkSJiL7v/K2wFd
JolcBHxZjd3xPpCQ25tyZcpSemqKxQWxMbQ1zKG1ZOXWQMY6DrjznfE0lPiYi3e1
gQN4lww05L5Tuv3HULNGUSeTdtkUuuiZGYfdMzSyFbOYeGSplK7bSRZPc8FJxziz
D+adry5TcKInPZCBZsj47/FGoMG1i1aV1/elYhLp6jI+2xkLWaLxlRVX9pLkvBVz
+yjBozuCbq1Lmj+oX+s0gBwyZ/49LT0c4zGcgoeIrs1X5KCeOB70Zd8+zdusx61r
Gd7mn6fexw/TLX0a0430jfzgDyL6uEiPuIvIfAReA25xNecpZokhUWsOMjGHhJ0l
+Fg1yc/QzHYXyYAjxbdZ7xaC6/Z4iFpMIJVpn/YYOrhkUf5T3ulAO7P8n1ff9tVg
2ffTzqEGMNdw5Ojf0p9MSCn46m4mtX4/Xh6w3YIgyTV07IL6+KL5BZSQuGj8/5Dn
sJzK/9C/WslFod8TxsJo+fyJ32OGpNAJsNTbk0A4gtm/a7z3InoLpUED2pxibhfg
DcSGA2mPlr83/i1iDO6gMtz1HHHAzUFwcmy3NQneNe3Y4D8pIATTzcuZ0FLugYes
9T8Rzxkcks3L73D8DIo+0zm2eFfhb9AdDebbmkRAHbDNm8uKiCWgIDAugjz7qNSd
khW3nH1RccBzn3CrXTNfaFbdGdi6CBz6cKZbhQVpg87PaE8k199HrJMucJkN45iY
sx3xQN1OOnyE6Er9oxrWSlDLnKSKHVEOs5NyabsPkdHKTSPbIlsWeuDRCcxTR3aK
jdYXXt24gnzCB4GJ0YkNw9rHig8RFgO+UP8dTIp5iOrKFo8A27BAedwSs+blX95l
wzD0bGCGW7YeKcKXWtOsH5YDkPUKjftfD8egEC/L3WTZeb2Kp+F4QqsK3urd/czm
qqu4sfH0NpHnxB6MJLANe4N6OZ6La3hU5DCKBomFCoM3DRTMyFBkzWfMWubruOH3
x1wDpCY9UfTyZfuFrgtynWWZ8dzLgWixN+rMzuV9WGnf21nu5SIyabxt8aXG3QTo
sO/9YGpFGgwyjVqG9gGlaI87jI0tebXMLJRA85p1FLCLsJbUquu4e55xvTJ/rdQg
zvOsbnK40OvjFgdlIsHlsqbvEhDJ98ctZ0HaATc0A0dY9LapUYOQ63X+FlYPWKEZ
hDmFvB90i+OJUD9KOdrJVxEVPhYbgQzqov4Jh2qhJzv/qo/A6kX4M01IZj8pFdw/
pVlCHUYij5Lf63M2KM/sI10Ot/7iF2S423y1C6Ra3ptaEXvphkcir60IV3r/zihe
1CGWVl6wDxdsHA5DiYMsrVomGfyFfZ8rtm+FZjgy31G2A3Nf1apMEleT+b/20ZZS
qQrBfqPZbSadB9VO4zVDdkuYYUm9fO8By3NfXe2rD4moJ4bASGweFmP85RjRug2T
/UXdIo2Nzf4zabV4fmna0K8KL2SSzod/ID2zb6lrTmby0dOnq2/kHcnGYeK+9fyT
0ny9no6cWY96cB2bVukxFagfWHPBuQC1s4Dm9c+k1+PBVyfgTkqmbc8tRlNR3cof
4jIMcYSjZabyci03fA4UJAcL59qgENj6pX9Y17E4sIQixd9kMTN1RNUTIJ+Krz28
vP10/Nw89/V2pq+dsOgI+24BEOp8kaiG7xyfxK8YAo9Pucb9h/ztA5Nx00Ol16Tp
YyIKFaIUdjGx0i9Ln52JQFd3d6hgruZvF1ayZanRHiY6BgHpS6RXcY2ruWIg0L9u
YXNopgfExsBxB1M93XGfL2XP8PM1pu1OmI3sXztR7xOeDKIhrJW9jZmHoA3y8GA9
0QaI3Yb3lhi92JnD5e7fOkcFt7I8vc0yBZrbw6tIk/6gTFOr32Vk/WbXs4gyBPMA
3TncU+2Etczow+NiGwyu3Un11FltaRfJQkIPePus/OAIfQbYbSCk6eoJXXjHHpbD
uXjzjNuBv8jBW7nlJ3meSWUaQrI9umTS2bdXv0ypK01v0N4ZoKCqbM03yPaK6fuA
SZ3Z26q6KqqSodhr6UzzkbroN3DtJUXI9p2eloGc89XFK8GsUk7R9jw8etPl4mGq
6NAIqc+iqT56uhYhIGpEQ9Zce9lCA9h1l5EgjVPjltmsLJBPNI6fKbPl9tr9Y+8Q
6B0fvR5FTbbp206nyqG4fIIVqPcRAZ5W3DONDLzC+xEcCl2M+kdXEwYNr426g8s9
84QGBs+4Wb+SK23Y+9bf4QOVyXk4tBariHEbckE0M4aO/RdNAywbGTAUezehznVt
CvOnJm9zwsZL7e2aWX+AbLuQ5n6cQPWeD6Ajt/9kXs4NOx4URqqJzVTCazGQzzL0
ClTbLtbaIvysOeFypDFhF7L9mHTFnRwwr2sqULgNKcgAtK6ULPM7RoqpAPbpiysn
Xz4QP0+4xLSpXdLLR6sHGLorJ2uugnF3XrUcFDEpqf5fKQlfJEOHYbYxUcRsS4Mn
LXmkyK0LL5y7NWXI23YYhnsM4v0DITFEkBvFmwNG2rPXUj0UDTP4Xo9XkJO6Hbxg
naW3Cz1uta35dnETvfhusoJXy7hz6LYxIPYc7w4QebTwEclxWILW4oagPPQOTV/1
aWJ7KMoakuMxT49CUP0ORDrs4TZWollxq7hOi+x1Wk8SzzVZZkGDEAGOempLgePB
LAMJgMmeJIIG/RCUpD+92+PedtYaAr8GhD/ii0Q/EBqCM+WkI/h7qJUHrPSWDLAF
eDi1ueZgGGcleInCjft1IlcuOoF9q/8cjfoVW6Zqk77iZIdzfl9Mol/VEHiDRjrU
YOD1j60mqNtMfRfHlOgGl6yfPcZmomVH3CgDCa9J7g+FVldeig9zUl6k0vsR7Zf2
a4eI7O+C0tGg8N+CugfIDhkSDz6H6TFbDKIYojGS5+AcfwI1eQbimbANxc9syXot
8FDFc56TxexNqo+Lkt5l8yRKK5LL2206KDC1tEXvZTZxvQJ/qYFve4TSXs0FDrFx
k0zlxqSN+8G583ZhC/0lGXOQEuMg0D5/y+cLY0H1+Qxd/gd28U51iACSYKrB9nas
hhgCdQU+JdkBMye1YXvKrcQaATYo5sbbsPXiOVnJpPd8TgYr3fPA+mKxbII1r4J+
dfyrsTx5GRY9VLpXKFw0RTor4j8F7zrjLgtti47BT5R/nsv53jIUNbzitJNzpNDc
hd5Ajy6rfvjq7thjAe9asz5xBFA4gV1T3YmkLs78BmDTZ3bsjHGS/UPcybFEaU22
0vhEXVQ0y2W1VRQ4cJeo9KLAiV1EkMgKhKqswmObhdFTzq3wMY9z92w7Y5H23dZo
ZeEZvd2yFi8GkX0m4MFoeZVAamhbTFCEdYRu2JLt9QW5CJ2wksmw97R0G8uwO9V3
CTYrlsw0FPYIy8kbalWLSjifW0wZ1ehIfAvA8Kebbw+K9g0M4cVReJJeNMMZece0
ZLU55Y0bFftBayjv2V7uS6bOLjJYKXYlfDDO6wwmcN/cdbOCEJvDU1ZjEo13CWLD
B4PWd7V4R/JMh73HSMecy324v5ytOFzj1A3s63beUVei+5EbarpNvyXgru5K8VOk
e+T89BnWS89o64kmd9vmPtOQj9C8P4Chad67diGA1xeAZk/0vKoqSNz2CkS2FIQZ
tYtRCPjXJKAaFPygFi7g4SZCw6VLmZP+AuBxD0y83YINhHPq4PSxLlSVwsLE5L31
aNlw9CeYY4yxnHcPtmwSY7iIhs9PDirAYGHYlU5rpOPyXikYqvXXuVVrq5abLjM4
V1dUkghVFr52R/HtG/WXvB8sNHjrZAnc7eR++Vv8/D3A4+7PS0XyyUdfnRDENdC/
g2qNVrodTNeMYYoa89fW2xPHm614Oj3M6+Uhzi1Z8O6kQWgeTy7MRV7c7IVCmMkr
8eKRpplp5nzR5Vo9f1vi1KICHr0UnozFdrLQLjn85WP22YCtSFdTxEwvTYsJXp1z
dXSgnpKdNW0NJ6RnFbY29cJw02HDwZEV5xkSdwQGiPKZZ3aC/GOj8Zbo+DY7fGlg
+2A294/jC/NESKQP/0uF0Kf3U/sLPtObUEb9lkf2nLE+pKpxKALdMe5tS3eRw1AF
ta75/xHD9d7a4YrvKHr5e4z19CuqEImV5RY2IQuR5tio5gUF2p6xF8tXpnuCcMOP
p/jDIOk9h8y7njYx8lpyWDslVha2btVnUXV/dGVtm01LQgoWVNLOejilgDY82IdL
fTzFQpqPZEVHRo1Hye/as8+/+D728CnpMguf+cYDZORsDeP2HksjK0zko6aFEpxk
umB+ZH93ZOMmS8GEwKYHzr0vH0ba4nLwFqcNo7kFTeXuyjSDsGxg5E6pbf9S26t2
SMirU8Z7tInfmUIqwrKd8LXysQFhHFbkSxt4XSxIon2AWVi8GrBb+An64jAUNWG4
sTlHUFn7IbrS/cFqMFY6J6HuB+zDDcjrkb1lcmt98iZRuY+lPMPkL3YaKRvuwTFR
iMtTSSM0qpjEn4h5SeQQkuubuPdMzUvf/FqYyD4BAa+c8K/RrrLMaj8vU3HjiM7T
Mi9LpKIEpWmIi747J6td6UQGWOqnY1Ss0GJ6wpAGMArs31IAG9SyzaS/OnYLANWz
e5MyP+FuzNR1bwTKM7SttXdoG7Po1KkpGZz1ILKIP25cRWwGqX7h7dddOR4tEnSB
/k317W7ctFk2IUHNtU8x6/devH3ucquMZqBDByfkvGPdF6+8fHuyrNR2mpJq0Hgl
RLYCNofEVgIK3TEUO1t3svddfS04gKg7GzSfFxMW15MHmWdH0su9A29HVPMZnz1a
cL4oL6TVmhPnoBNBql2BDAqfjuS+8d35iDeK1fZZUgjG0MLA8xsA4wojMyNSoMZn
DnNTaYO29A51bVIt/yHqTAnl818neCeFA2zgB01odJSBqC2bQ2VXIfVzcxpRMagS
OxeAEtuBcTOtkK63Ilm8WxG/eruZXPE+Nnflv5a9P+pb36FLUY7IYPmq0gu0dgCZ
b0SvRqKvYYRJUEkmW0a3rq5di9sYvPjeYafouMCQeGssgwQuVhfZahSYlyjl29A9
jH/bvvaS7jvUhdx3PUrutYVN/CceYMY6HLaOX5a+0/KZZSrnvzGROvH0O+w1PJif
HnsXj5dZSvY9Rx187hx3vFa+VMvWnvGlhBS/l/c+OF03+q6f+0P7lRt3vfANgg5X
clSrM0Ip550MRVBA4CWqyoVm96MjGQ5YEhJYJ6bRHUgazsfWNDRIu2d0emV+Y5yd
UIRkXfU2D5s5zdN1wpXWIATwCHa+cs0Yifh5p9xiyv47FE65rRa/uPNFYMP6jwKb
NB32U++6kVMZRZ7agSpmQfhqLYN5ZZI3NtYHZJqOnSoESy07X9D7I8Ln7bWeNPf+
BvuLY4w7smySrof+tQ1Mjvna/T4nveGOc70dEuGs9K5g+39jHxxFewosvJtYZReS
JMlVrD8nwbM7D9nSbBoAq8OkCnA88BiCbOTxxtHpXJao7tsNrgBVk3Oov5ntHmQu
JRhNkEuhGmETi1nHd5PcF4TTyPtmo7TqdGD6Zn0alhz3QaX+BCEIY0sKXrDpwCJE
v75FsrRyB/usG4JFKaxiNQbbxik3uIGl9cIo07/xBTTNlNVs9UArCgu3OKmgdoU7
T82cVvOI+hs0LaODolOdOhjUTbPWnupO5SJE9GXzlP1V0BBbx8DsUsJyOcOVecQB
YEUXmGQjeqQH0IHUkwybi4Z3/yc1G66SfoLlQ58SJ/SoAK3Eob8RykDTPhOm5PvS
6/BVbAf7Txpq9Qj4ZaAxKB+QB7R7fRAaj15rA3R8MUeY7tJyS+rAWpnonbgnLaSm
/MLxzMF5kfoKcy3G+tfTWx2xv3PWZZWvZg/PJWwJKOb17Y2YeEITEj+S5y/zvYmF
Q1ZycqvXk1XTVmhUct+84lM7bsqrYJWHs/weQichEzhdmLO7FpLdTnKFqokPm3Zd
OVz3eGuS07qEOrG+KsVQj3npux5KmUjCvn/DYwOGssibBui4TUsA1PCgiOloojI0
IfIIGJYJR++J82f0WO3KkKc33ZCBjkldOQlLIGXfbYhnAKMHGbvRiBz0cfWX5oRM
/NYdbj0oA5fpA5kTMPSc/YMktRF1bXeC6MhAF3MuKxUoA0vWOV3IhG3PdBcBs7Mm
TfXDMBHvhgymQpkXrEoZ67nmUnZplq5V5NjhTEy92WRB9V9UL7PdKTNkO/6J7giY
eTZJk1yjinXJSNwUek26p/L0eagXjpHtMl0AhZEIN2wV/b3ndag7Mja5h7eSgpD8
K6T8JpvdXNZJFuZao9Ly0VWIqWn4dfALFhldPxxueZ6MuVg1wjZXejdyuS4839u1
FCQQwpa/1KA0/JdKFA/kWDDWeabeEKXbg7KxajLmAb+ls2SWcpAP1PfEBxwSoZQ+
s33mWENKPj0a4DK9gs3aQJg4GFd59mDpeOH0RDjT10WhzMCqfud0uaL7jQWE1lYb
g1SBGF+UoZQKh/3xRhl5AN++Jj1CxvUUJNGExlRCk9QFPAeizwt+EGK4/MdyhQQ2
B4v3xxuGLhYoTaKrvJOtsPH830xs6LAPi65jjM2b+LvqpoFqnXhDmdKYJv0e4uC3
sEJ2A/MMH//wdVsoKXJuVl8e5WhURQr2IjgG9tBx3i4CUW1jpda/jqH01d1cG541
hxqzzVJu5ZKyEXuvrw8MZMtt0F9nCUOL2MYQ5mHT4EmBlRQvD4sHPRzzsmi3/stQ
M0ulyftXmSYZ0977PAQe7fbRcjV8otVx1CfBdcIOkvRwwkfYYcLEhf2g+W+BbwNF
4isQffuFXk+mzLAB/ibBXllh0z1ggbWcyYtWE8E2tbGxlRinHM1dATAksqa2hVYU
rOcTukHyCVdtDw5WnQBTpRq6Wi5OViNp4TFxookjZ8oP7Fnfyapojbh8X6gKQfD1
jyivjXhESwbe1jsRtlIvTamZRTQiJAO+Wx7X8KJl0Q4tY3qTPkZWoR/1JJ2PCfky
3YKrA7vBIiRIuzTXofGg7OvVqnSKyHzyW6J+C7eFQ5vKVbxWqbvnJOOnbB7CFiqZ
Kj4NqiFXanjf+ilcCrK+ohbAT74IKdPjV8HJ/4knQZUCYHp0ruGwFHRM1tkNB7PX
1/gQ3qVNAaOd8M/tv/lIjJlBuyY0kWTpi98GghBE1woKRfGZtYsBmVucQiYWqWqm
x95HTscFiBBw9+PQIhrGlwM2Q2NiK4CxtLDhP08EZCFLRDpYqLLrfJKoPXN1ypTN
50Y7uVvU+no/L7LmXrVRLk/bBhoWq7ZwyJ1kaYbtgcrFZfcaSEVeOKJgjxykVMf0
K8S1I4YqBNaywe25iQi/6o5OumsEaWjXFrZ48pB5q8yPbkVnx2qx3fJvfHA7/p4v
dUiK6tgXupoBeKFdbJbZYJUjCnnYdON1ilXntmMxOSZ7IHufl4VwiESelKo+SO4C
TiKsoMBUTUNlGA8XLYmUR90zXeSQ8zktC4BJqUVs8cASIyUeE45py7IEFh4bhB77
z8wIq5aTZLB9hEK5ViOqQvu8jmA0bRwR+t4p8HbuUimVLX/Fd7fM+Bf5ffUOld3f
b+0VzE4iKsvb+Nszlpk4aVL1eqfLoBiPVTh5j25Q6G0tB+VlKhvhP9DlG+mTGX4E
NxwnA6ofYVbsa2WntDKsmpx+nvCD6PZGIBzMPCTvpqiWPpo36rzEObetegNnn71E
6GeSiK9qPI1ABtPfYi7fBwWMlW8+5lWgfC+2eR1Vg8s29dJg5ydjqnU7R6qBfNQf
Es6f+Vrkyp6LnOhg9tWnJrdW9dQ/ipNf/d9lfQYB7CnSFWTX9WAVTzdBhXv2oGPq
Xntffl9+jFX4FegwYJ4aYZmL0yIwySLGBg9/n6OsoilASUuITmQnTwtpzk4Ug6b3
8nwntlkX30j2yFTVMfuiHnQeW0mxuiovCze1OdDB0JobRmmGI4dsPtrrQEgjPaJX
mx+cExITlM5j3gmoN6FtR7FtiHOZNRPBOC5D6ePCXjJDrqwg71xqKZnfjngorfPk
exMya8Y1y+n8IFnR93oEzbBwZgyRpRAD7PgH6wjiYQIyReb4bB5njaOG16509UXm
XJdF6+5gSb2uOCnE7R0cSdo8rcq0ixnlrdAb2I6lKmyoy4XwEoCo6Kuj8HoOO4Z/
7F+V8cFaDLonTct8ulJWFPfx9fxAdcRkM6JEIyOtudarRTH3PldiI7i54+ZTWgkv
MhegdmaIftdZyeqf466sC9pKEWLJ8Ak7ZtH+l39ezQqqOy3s9L9omVqDMIBmPIZF
iNxV9/KBpaUoqL3RgwfD1+TeNrW5hZ7FbyeG6eAeHc2DkblveBQvZL2He7DrYgQ4
3l2dWvzGzY4u2chiYGcucQKg8xpV2MXzbdfXTgweNVqKsUGDvOChPegHQXBtvtBH
2AhkBaTIF3L/M9PKhJoifDThta7Tw/7dyBz3jlJSNDyAtr9nebqfd9f3tMn2BLKp
RktHKfxZeun0PiPs+PuUDGWWTy4D4abHDwybDL0rpZZ2NC12xIUvMapDtsZ98I2q
gjjI/Aid+mj8MdcbU96m3G1Dg3TuRuIcTBZyfve7DUWKbuxsDrtiMypkQ7AkspuM
2KBrqEYb8kUDHPgIEMx9ihIA3adOKTudbv6aUmKrvDznYh/8LuQirZYfa1a+BdUt
HIMe3m6vT1AAVFQz8SKvRauu851ZsfsXv3o2Me6zgGq5QreTI+Jy9wuxK7KvSOAl
pRR86AU4pxMBjG8Ca+KHYd/yc1H05j2uzwdZTF1gcz1xgPHqnFFLh+Mv8dbvpYGI
Bij3PARB/iUf+XNDbaRLYeSePshOPjS2zn46YMqAqaN4g2wv+nU+7tOuESx0p5wX
X73P7gMaRPaSc2KMJY1cE6lHU3Tl+hrvIfogHVcM2C2q616jmTL3Q4FQcl5GfCjP
Y3hVEigGiiGn5F0+zrLfPNtqjXvCmoKGRjhUmvaCN6aJgSoUt3HzIJdFbH4VXZU2
md3r/Hrz1WwNSL8VYc1QPS+s22uO44AumMjmChuWZT57wotkxhbte8/OLbU+DNdv
OQbEQwR3SYzGy2yuXzQqmqrlDUGINPW6MM0NvMuZgrlG3T+ndRfCpFci5nrPzmTF
x66pccjhQji/szAQcv322V45ShywPy/SaTZCnsXiwbVK40R7DEJ++/vO+ZPBFljc
aTMZ+ED1GlCsgjgNEnK3H50pAwHbq0bySQfzKCMIqG5poGGdMKoDHK2wB6WpUSek
Y9pyWpDNkSCMgqO3f0ctcevgBOuWlVGvQvr02VLkZAMv2qe0j+VecoOOfQ9CVy++
2NOXZR3h6ZYDLwHMkHLxakV5YX7Pr11Hqk6YXEULbna/0NIXb5+65F7O62oP2dw4
78P2Wr/z4kvaxvWyx/DpT5RhgexsDmtf+CV4jKeAVMq6wA0HJb3goQql4i4GdpmM
k8iZkGwHsj1WJ6jiswTAp4q5BDKeDhoJZZdEwPgUeHGo0zXN1Gbs5Kyx3Fmywcoh
cGgiSNFhnexVnLaKeclDS0yJf6O9GrFiI5eT29mBCglv9uoVFFI3P2xYOCM0Klp2
8dlMcClFSjL7vgdOvW0nIWj8/ym3gPUTJMzwsgm/bXOSAbhM/cgEZqLQ9zs0znSe
6NnSMbtXjVrH12sBDUPIu6CGJETyH4BR0RBV/GAcDFvAeBArNuCR7r4KeeRLRN+W
Muq/mNhtJWQeA+uvo9xOycBr9XsK+a9c5//NNt0TJseViOmVB+Iq5jPuHcm7Xrpv
ZbeHjcFS+018RsipUitApBKvgw3wSqtFSNRE5Hu3vZdNduvOJ2Xt/3JXbIBOeXjD
By2GmCQtdRlAY0cwSISfEmpKceVc68zngn9BmvtuC4d++HhdQPe7K9NiqZLWDAUR
2WjLtBInzGAW//ToeegIm73vniKkB5WlS4GpN01rGpi1xw38Ki3GfT1/kp9lh3Gu
gk/asOKPE8n49oL5u9TPNzT7mAlSTke0Nva1BCBFfFEV0RrzbiY/6VFm5qStxq37
JjDpdaGnPxZ4wDugcFh2JoipMSPVojNaE/diFiw091x1RV87gkjGeUUyLi79Olrw
vZX3jMaFh4mOQYt5kOxVOsTo6yVa9SFUIbnjlgr+BKfh/2XU9AJ61M995DrqTxIS
jJj51uOQGZ8uAli4jS/9/V10ntjloVco7kQXDKX5Fk9d3dRo1NcWWnkP9oKhw7a4
hbwkQdEJJGbiJhvS+CTBOgpfJcRqS3T/2yXIWel218A+vAX0TXVVOhCG7VjCvsFj
2OjYMjEXCt94eohzGrujuZGSk8Bcc19VkYZuMfeYc+JlfJSvVLmMs988S0sd10gW
d9EczPvldG8kDCxj+F3Er8Xvfkm9ox5bRIT7609QBFNqlJP92howeebEavk/fYT1
v7uARv/nCVoJ71ztoMtd1tqAQ5VcoG+YSrn1+lzTNPpvmB9nE7730Au5A2OZKJB0
DBolGaMw5//iZiXFM6LD1ahQpisQ2cRS1Qr8jDSSM8HRWR4Pbn3N6J1JoazZgMlq
tv4KLE6kHO9007ViBHCUXruz+AFOCXOCOZGY2Jrb7ilEgV0UhwmfljRqlyt7vd6W
ESruRPy/Q1Hy4jOD6T1K/O3CwSnkglVC8JQyVAyKz/AF2zSUNFdZkHzQ3oDVGhZ1
TlT0lEQ6a2lbcZ8dpW4TYKvCPsjs6xqkMqhicDkJE9gCOBm0sFEsSUvCVCX+L+h1
tdcjgdIe5Thwkv/7nYDVzM0tzZGykENRzXA/xLSzSIf1qzKoR9A+fL0NuBVV1NPr
f9TqLQ8utzTVxLQQmOrr6jLc6Lu87VgRUIx1r/ry3957zV4IqDHHjqRTReemvmt8
XkZJP9YrPaguGdzejmHJ1jobd9fe7+4LVkpipI25TkRhj0Di6fH3BKL6ne4ZsTXB
PhaRSGWEkwE4O33xjJIXEjg6prHAgM5tOqKk8xk16/YyF7jer10jyv3AGOPz2mvj
YMyKk/nOPt4tQujLE4IC2ga/ozOB63oChEyNigEPja5PqaIxW8UjR9GvurVkJ+IJ
Fn3du9LZ2oisZoSGh6+7+Qkz1/Tu+n7NHzgbYHlc/zrk+gWEQtIZvGTY8N8lta7e
f3keCZXlru6wPgjN9ZSR0sQV84iWWZFQcyPHjYcoc/rPBNT9mliazUAAAnQDv3tq
uoly+eX437v98tUy/kHqus6XrkEPbjQv0Qq8uXp/AzikJqpA7hP4s3EdYXzAqh+x
jlZ73o11TTyHNkwhTsBtbwks+IGATzowBHyknoKYM342qnu7G532rWzsbFXPnV/s
Gn9RaXksHOU2W2499JeTBLL5ZoAbNt78/5pZZFiO0e2LBGSc/mAZcGmvALL1oNcx
3o5zqvDFAymemAv7kztp3a3bUPdxmfaaVTCKRogpJsFovkNthPb/TxYlg010XDmd
Yzq61CrxFZkNfQaYNi7I4y9XFPULpQj26t9oXRik46gNT47rR45y57sQLeCP3Gvc
drNrZRoLlskHusCqYYKDG3BhBgbTwfSPcW6z1HMRKj7lDzOR+ZUgwmTT289Akluo
iYDo5UuPtaGJO920DhYi46J3x/zGnP/TvethlIA2CreWbt8kMdRN4mY+aXi12301
Tytv5xGjsbL06GXjfREz92low+bQ2NwSPwxIqVxvGe838ADRQYody4cE3B0qZIZR
At3PNWTQUDIZ+Vnym5glMtAAgDKGO3YKyNH5oHGDrLCA57r0AiMWX23V/Beid7JM
EjtreFdRAcmLFZDIZQQtb/7YcH+sLy/1UQoZT/U915Hk+/scLrNlT1TW5msOI9qR
0KcK2YmmRcK0BIwVyXv1ig7X5YhaWq40s9WOyDTdgNt1t/4RULie1IA6lK4R2PSY
ihWkCpnoGfJfyBDtCTjETUHJE5PIGmbyAZD9iW8jahn8jRd77OTvuLufugI5t6US
XAhN8HsCkpxsO0S2nthegWmPz7rjGy5pCP7y09MmxydDbnvHpyzE4+hzQoqqYFtG
ROHSAaXiMaGQBkjkfEXDKeD/tRUZFC+BUebt0ufUSKGoqJzLRzrIsmRa2mhpxk1Z
irRmIXwt+DBP4d20IFsRnm6muemK+kaRIg7/KK3EFwTUIzwOXeyclgchx7ckrBLV
R/mI630HPnV77v6SzCsy0I9kEbJQrLUWWgl+h3oe81d+uuvQl4agkzK2vWJu3qwb
66b8gsyzHfCnku2fV5xq2Qv8kWlg2yFQhCZY1WnraKxJt5wP+gbWp7L6y7DnxmY3
2VEG9+8Abbsr2zcKV47njiOzElweQIyUR/guu0RRdoT9jGemafh05/eD33t70U+W
t+cMobJXho7egHalAp/ibmwmGv/kYdbDsxaqsskHqW+didgrTnQKAx7YPJgQICMA
STrtkVBOw40JzZXbhm+AwRI3zLS/bdrEGCqlZHp0YDG+pk0DWWYBSgLfX9w3LWst
jF1pX52QLpHKi2kgG2s3dptZqYkD+DipRwM/3eQMom/qAoz4Z7G3vD4HzHv7kVu2
bHehceQehkpu9dIsaFaQCDqSXaeLbY7eBpwYFF3svf9LuKw3ANI1epeAFwoDKVns
CIy+rajpC+hkkuQ3ZQnYZUrYOanFPdfB5ciJAalJKPeKjsGzD4URgyGrTEwXkRHU
oI5oh3BaX9YXPLiePkKrOIOQg6AcHItOyDF95YNe0pYqLwJby1ao7Esrtv4h2ZpF
eR2a8G/bHW4se0VYMy3X0Hhly40tY1gwBNjSI5M4Q1e+TWt0HE2GqqUxDiC6k1Sr
z1K+waBhbJURW20eJrbzf/zDy0uQlsY0vZc/ufIj2J8Gf4Fs2cRo9LkmK2n80vto
fKMfQu+dKR0zU86pu7qJziU8KHsgbE7CKhMssY2rbL8J699onu8ld6x1ucVIvnqy
Bd2uGFpF/rHfuqEeR1ZSd7HaMTUafug4wqALhlu31dj1ON8DbBNEDUQXBGDXHgMJ
s0g4hq9ITbQeA+IWpSSK5OPXk5J7ChjDtyEC/BdP4WxdiiTcJt8nFma31t+B47G3
6EhR8GMq2ro/5+mg1YSVLLuL0rgKI4rN3R6EWZCOMHyvKbWdflGI91xXQj1BaRCQ
YdwyBeE9C/otUwrr+G5A6CbTMjiXx1GJ41CwHBjcpxsc72L+1JphCqjDS9ZznafJ
CNi1ijEE3lHY9CeNqFxwCS510wGC+f1aZzfkbQR5TDEwk0WPS392qOX7PH0t0JuE
ljTkLeVchH6n8HTXJ65K2ZpH7SSiYkJvs7EuDZO5hHT2xHwy4LzNnHgEgaCRS5qL
bNSXnjUiIGXnDoEy+f7vKhn8gMjPJVNWjAq2AmL4ZvrSe9MZ46TNsX+SkkJhc1rq
9gZ7c2aj/JtiN74Dkz1OhAQNG2gjHiwh/knD5w6dNhqoKNb/efgqrPP8lcKEgt0c
1EhLEQ9g4Y1HZ2WigEoAIR3sO1WjOzLV/PNplU+s7EtkDL9uuP7/tvMR7Bqq2+F5
V4baOiiqlHaXCAOKXhZrn5cMWQeaUGY2myZV+u7Nw4143mcjIJy7tJIxBqg8pSX2
O4bdo5Iy+iTOhHCAlz0aSeLMzptFnxuDZvFrdQgCU6kMvrLJ2NvEpRFtsqyGpk9p
gwoKHgyySDQwp6fb0v5lTAqOVJjpYQuxmdLIKGE6OIE1rePZSH724LR3mk2C9xxr
mLWnF/9G7gsisq4HP/wOpe9U+f6hvDb7Bckco9ADGDZd4Oueleq80clXU85eQtCT
wKC542/tsbk7jeLSE4OpAvOAeK2h3WXwLNzdvj6Kiq/E+6cuVCU2Kkhdf5OH8RYj
jcqQFOuqgD0e8kItA1uoMwJ4NAXSeERk+dYN2ysv9WVFczotbn6l2kzxpUZ/xXZk
5Z4Fv8TndNYT4n5iOcQECfosKOOujHrUq1JitELs2iNAUjB0317yULtSFs884ySC
BXeHKbwXcOo2NBCJKppFf9oBjMxix3uuvb04M8sKVbRADm/vP417ljY705PnDTTO
Ag5EkErUD39eI+hkUT8AX4xfPSr4Pma6YGnYrdRl8wnTuy7FjEjwuJLXld4NXbck
10pSGUgR7jstXBF5BJSCRm4Fh72DYw2Ja0EuTE74QnLOgRhpGFQL9GV84L1K4pnE
u9uEYkRbY605w2QdGrqe8/QYmoajYhtISXKuioL2b2zfmR40iyVPdTM0pAgUUyl1
6f6lS9m3uQkMBmXtQNdD/cmWb8c3wvEEsklbKUw3+61C1waUkOaYUNijCaPDRU8l
f5LnALjKITDzxf6KHwnKpsDdOl+TiIVPSgggVwFqyYjUJmfSvTcmuFu1CBu1vTBn
MpiPeS6JmLAsHI7nEmBI5f2S9ZdHRU7zY8QAzrUBWvynZD3pgb3gUqSmVja97XTK
w6msmfiyicx3HgwUMWnbG6m0R11yhQ9iPEzXoz8ZnOJSDaGtGw53wKvtbiZdozC3
U8XHdklfXs2wHOzfdhQ1+IKhL2Tpu5Lxb2y6Pq2q064WWiklfZNH1+qi6utn/Szn
NWsK0sa1FYjToIxeqyWFfuveemyacZBs+v4r0cdm0zLd/DdaqhwLizv648AwG+Zo
KpWbuI13qf+hpRLOfBuukW6ab5c6Jo2l4B5vg2fxwgFxqRwq/JLYr115lRZCM/qx
//MGhBuO2eVerra/1JViVT9/y+KrUHLs6fiE50uTu0MIfL0nj8YGR9IHosFG4Uir
KQa8sX+ZR8JuECCTdRenvzVQY5/MQ/eUTiv4QeqIgjwajg8mVbb1Iqeajk76MG9m
rEsorJ8tIhTFro+0ka6UJvX1Nj7gMMUznnfNqLY0W2FWDUc2tiM4bbSNQtK0zFa3
jOQkM5ukYIfShr2NBlz+HGJRZeeaRy02E7WJ2ly9EeCx8suZc3EdrLkTriOOTSbX
S5iItChp3Lhq4Cq24OVDICjUr5c0iPJbFoaXQn0dVd9lJ1H4sYwLNoATJHohT0mB
8aA+c43VEwLL13BXkvCy3QmuTSObT8AK5f8G/5txelP3MnR7NRY4p0gU+ygS5HzN
nShEwEUwZJvRf2ZFNZ0cgtiZiAhR8Rpzfyt9FRWmofF+m9Qj6hzXPdXmz4DQ8oHo
q6tmDIl/YHjrH28AzK9c3qZobDu2Nr8+SUXfNqX4vuHP1zNFQt+qyv5Lxxiui/yD
lr5DDpX+j/upY+kpw7BUqmFRSo77CiXkaVYOaxZA+PPShJaOS7XPSkfdcSidoHiJ
kETjxLYY82Ee17WosyPvUaoK6k4fNEEadaLk6fDI0RgG9p67bVUsNtWGRCIqvZMi
f+SMUqEViS9ATIpg/Wy1TOBlBDIoYkNe9JV5mHer1nC7UhPIckFUsN+O/QKMMoEs
PGh9yxiyz9FU+tGlcBrrKuiE2zVVPVW/iDBy5oTaDURzl3x32Ipa93mRRYvdbQ+W
VvQ70c+ZEBm/ZmiiJhRc4A/Z88t11aZOeX3JYR8ap7+IXQkDVcuTpjEHdA9mOlN/
At0nJufcHt7Jnh+ZBFETlnamKDeuo8OsKP7bHyEjNQp8yqUXpUP/579OJ9CCEj9u
B18porKfOQVsLgLY7MAzgvwUjs+kYLVNE7Qfx8aUgAMKcMeDCYvhcxehlIkYLMVB
GDVQm41bWPBQ0eGChFH0riVt29YQ+ooza5ipXOFI1rkCb0Q/pNTYRkOssb/ua3y+
/pS+vDbA1UiSSZOx7ptvnMdQOZrMmwWxMcOke0Pa5EVcsrPiMInGhAObqCF8zoyi
dvh5bl/uxXFrpZavIeAFX8rCNXaSEfR/CIHrieX1cC0UD9iwG8WsCaNS8wVYepps
Xi5qF5FEaGRw9tfb8ynPh3LFfUAzBbEqhjPDgCOO0D1VX1phKRTaAq1lQJ5mhCrX
seA3MpBcJknirL+QE3FnLOsazGFqv4FTg4AfMGTyd5mVgW7ExfXxn1l1eHQKYoir
kYjuJrKKBkwrN7uYLfJRfc9yoBFQDe+OIb5b/TjyGOZIoh4Yi2HHnhLQmdMKyv8K
f6cpDQUQIaywLWVLAA+ZBSDSvb9YDEwpI3pkglSWEo0/4xlMIcpnwxJ7gU3D11Hx
K/dJ4gpi9VqJzcVsM6YWEJKDi0ZYEjKZf0V9u2lMHGXT+Nzufoz1TJFeQs3l1d1P
+qew4LN7DYgpplXVAl3U/Z5ILrY3/6DnyGmTed8p/K/vuxxyHbw/wPR1Im/iLU+Y
qHIS4FDL7X8n1AZ3S93ZHF4VRv6z45CvM2JimzD01CHO4PxUXdvuagjOT7rD3JsW
ZPtxasJE8UwRhtwRhysW43crHpcbueET5lgP+EyF1128yN9YeCCkfytVU6kd2e08
kgH5OMe2ewtTCDBWvC5PFQPcA4J84DTXq6CO1hW21L6AEdk9YBVrLbyvh6gTD9W0
U1V432Zg2bsb9eqUSfPVKl5KxzND+3K+XTvPfeiAo+SREKM1/n/ntsRT8Ntko11L
uXjFEQ8AuPBTu0oNozqWnRXdYLhIQiAQwF5WQUs0Pn40v2l4Eh+OYVU1yh+ERmA5
6zkeZ7GjmyTUOtMbHZpFpNRIc5fuEPp2eXP3C0nr7OQmtNE0Er5VnKQaZ5Gfw71M
hZV6NpFkWXOx6/wNRYoGMCiaYJrlfX+5gBkbFop7YEXGUCPFF6vI514iNK46n4VS
SD8elIsFEjN7xkbgpSYvVBc3BcnbFFhuZh9G9Atnxuk+MBBnYc3w5/pHfIZ6RQFc
QEDn69XhjAiucyjEkr23cAKp48GB9SpLlDAnVSgygjAxxQmCADJnHq04tXc57urx
IcDpP8pwTxWaREaTxMLEZAHI28GYyf8WOOuXpKgaYOZISyCVv1WKciqOLJhilUkK
cUqzWsBg7AxALrQMWKyXBHzaFKpNhH9ScvBygq5y4UZaBDYhgQNsyr40/LD0u5kA
uYAeEQ8u5a35BOGogwJLPBaZmbdtEF7zSVUzr9nyy97NoHENHG+w2E4MJTXEpVW/
pWoh+o5qMsj4sPVXpNZG2ECK3voCl8MZjgQMwGJXZsbsUnA0Lw0jFp5BHBoWbyGO
f+zGcARgDojbesD0lOBW7d/BE3eL9gj838jhe15NdZfexkOHNu7NHlXe/PAvtyNv
X7yao595nfC4kPoTDyp6LSLKK1qFB2VLf7GgH4b2wyOjPXJDxxa413BvtHiWcyIW
sXhpzW/dv03b89t2HJLkVtjZJGYGkQ3JPpPE9M1b5a07Z1byLvzTw54XhaXTANeG
G9g/64ioDxiqjfbMSeHDxdO1CaWxR+ukanqChCaewc7H4x1ZtH13v3A1Uv4i+C7q
9EqH3NaZuP95DB6gLFNpe58c+6egFr8fBsqkYIwJUsqyWHcqxypUyyEXQ3D82Vqd
Ev+kshM3s/3UY64/5E81o2GfsMQG61HkJH0SMxE+cCbi7645e6t7/Fo0qiE3nMQs
hmpzvHPRXtSEp9G2MRYlsXHp6A2nIboNWld1ZPlGkCuKcZ9XabjSwhADMvZ2aJR+
ux+vdlA8SmZsbEXfQRDYXmGxwsLykxv4pB/efn8IMsX+xCjJdAaJhwrGEJfT8dcX
wDO6OzfK1zzidlvy8qgAlGZVlfJkcjNcQdcCiFjLfIPQsDFGW5lv3djNEmDhrDm+
KeWBaQvTMHoNPAlcOOz6Iqf+xlkD6uSEZ2m6WjXsT44KP5qxCRfFj5w/wO8buhV4
1NujMKI9cZKgMjy8e9lUIiAhvpY6XqBRimhuJbGgx5jNDC4FimSPJaXYEpzE589d
j0OkyH5HPjLHCpsB/5ftsXsViW01BDvDkt6K+8b+12uyXZMxDPBLfNVCzATdSdsS
e1LWbTf0cGnlP7wwQGRUE63TEYVn6Caay0sU3Ul3ezkCrwXs893PK0Dr9EXWA/mC
/M68J18YshzShcnKr7WlQ9NepRCKI5PX/FQQl2Bd9Ahok+gHgjgptdI8cqpyJgEm
qzxE4MJM1qNt+h0pHvTC3r90rQvSJnb4aKLYek+bPaBAympinOLywsm1hLRRhSEz
oa2vcLFwPKvBk7mFfd4ghT8SRYM6Weq9tByFu69h76Gx/+Je6U9zzcji3zEChnI9
fv6cfzrYK4IzdlcLlbXceYFA2KzrJj0GlStV6ZToJOkAblb1j/V6YbNpB/RgMbdG
OS3TkHbsjyLV6qFgOCmzbKE5dX7W12J0++ChNxm9x42D+TqIk1fHZNJ0YiLH2xxE
1yzSktiRDkxLEIr1X6Rod3+Qza3Oi1VrA92miH8YJGmSNAC6ZwiDVFzrd5RM3GNS
OJOqtbkJIOfVNFfchOy+cI5S+d+Kf93w6WihXuGaDj2RTHK1wXtBQWQrkhTSlYJP
1LixlFtMkjMghTp7lph/r7o9pPlmjjAqL7sBYQG3GPUPjyraWsyxgrjKUcNvJQtj
Cogwpb4Qum3i8Qg9DE1Iq3nKZkNZJ1bFvxKEqlS37JcEoFklg5bbgk7suFR6tlv9
W6j3X+5pMLR+VONGqyHmvBBBdlnoBZFymbCqenvGfhQNLLEOBHK9xGCCynyDFvGK
W3DivVupjCdJSCp/JwqvYcpNmh5FAgA1gKmow+iMpWUGEuXpIUFKHUgCESwodKj8
xpjCMMygbk3+6LWAs44lJg7GOp3HKoiHNAart5qdJTe2oxcPQyZ+qXXpjpY2njxk
FhmQHzXz1y4Nb2LAeGCsq7f/DtFBtDBeIz6YWuV9vUUmleq/CGJ209/69fGesfwA
i7N8Pc+SufhOGWtH/CqpYY/Kygv1dSoOd8+eLXZtodWB7g808+eZ/GjJSMwxfPg0
OLp7eGn1Hf7tbr25oMoiq1wF2N8oon7XVNJ6QFhoQPJQvhwuAx2yL/qsiX0Q8vca
1HNCt3f3tel2sWV/IKKl+5RmQnA+7140CvaJgCODu2I47vbeiOrTYWLiOVFcmt6W
17bDXPSYwBjwI3zRCYt7jy7GNAlRMZPiokQgl9bFGxTcUsdCvtCNaZu2BGBn8gCJ
4XXwVJ0lqr4j1Amq15q/b74hXQaLaBza8B2nGKMSXA4wSduDk5AasPWCVwi4ZnCQ
h4Aff5QuhvTanK7DghoYZv/q9Ul1xhW6v51hgtgFzLWuuWAZpVJL5OneO6MWjcK7
zIwRjO1OYqbOkDXtKGYDAm74DdQczpyFE+kJxadHBAFT0eNmG1iukRtGlx87mJSA
pU6Dyu9lbH3A8KBSAwykSoeKtWB4wKrR51igXtTpPqvDpnjejgG5FqQn46nfJnUj
czOcXXDBH8BhrlJsGAX3rTaF/ZZE+9bYlWlm7Hq8qfqdlVri45SHOAc/w8xw4EGh
S12Q8b3iPMTJgh8RvoDOOpuCPKBE8KmSKAip6eVS8/HoFsYqOul6+G7PTO4+Exxr
LlUONZXS3K5D0UhJTOEIhLfBxXdSRa5HmVtZce2JCaHLdj2pgs2b8KuiVF8vth3l
TuWWhbr5F8uRy5WQtjT8A+vH2AwbQoASbsCm2SuYaPtsJjEW3j46ohtuYzZIqF3b
kDdOglJSuJ3vXVFvGU8AavsgwgW6BLMg0C0j0TJ6QAXya+EWUFr3gjffPdOXnqWE
WpgtJagY6Sfz+r30IhEqd4bvqMogl0HWPZtMTuazPFDfXFENsjfzA03mmm5tabT0
ViB6Hp43YZXFtDbPEiGeKOWkf1ZiZSrM1Su6oWhZ8tShsrzMMpRur53ckjP1g2ah
CpKhixMTUN7IooaVbAHD//uC3naFAsqZubLmC68eZc0eg4ZjXe84A4Z4JmwuYiR/
GLPFMz9UoU0svbsbowul3uWoL3RIyp7qryKZ5Z3Pdv0dKEYROJp7hi95uCoRLBJI
S84ZkWmnx9TGkwVX1RqFs5T8UKEJ3y19lBuDTt+WzyS3bTF4K7NOq039HICUHHRN
KwxSLyevmpwi5dAASufmRheiTzwMgYxrlfpyuwviR1RynKjk6KVPE1WWrz6g/C+r
vaQWB8tmbImlT7A4f6W3rkBdxYE5xN9e38W4sYbpgqVW28eBDvEQ9Be7XI/3TNyl
x6H/+cbuDFSrVTZBgl9VcUrWGSS/Wlo3/Xdu6IFxuJ1d5SSJ4lATEp6yjpboZMdY
i9Z2phAHHw7SoEZJE5HnfaUy5djY45augFWNJ5ASWCJLmrkARXiV30prE+Jt0d02
dfTAG3BYtcw2xP9D7krBWYHMWOcaB808yvvEKgofkFlh5KY3fIzTiSr/qLwEpgPT
mEy2t2y0hRpOsx4Y2SDpHimqL1FbagVGOemur9bD9rwi5t1fvw2a61l/0+2Pf5bb
rv7z5iu1FrRwdCAZlj9szBZNZAoKtC+KeWW+5H/MG814qK10DjLAsf/WlSkyjYO+
fV8ucToW2NaT4gIVsPu/SzzvtnTXAUbj5hOxJffNnwduyPJOUt5LqAFTpZlYFnE+
KxLzmusNUt88trjPP7cHtDbB129ntykWQbnO0WpmIP8xiM4tq2aqvuP+DplJTIVf
BCkVSOdaAmgNbFer0fuL67qUFYCeZj3f5Ws7yg9At0Mh7QEYRJB6xycoPvneK7HW
/okYPef1oIPtFaUzj59Ab3EmtXEcLxbqvtrPtEpH1G26POJJvyTkI+WRHaO5jnOP
usBNIqL6urzR4DE8AAw1qe35KBziZaUDJyy650/FxFzDB2PfyBJX3JR/iAMwFizO
ZVpGn6niApJGV8nR9rWRJZdUzsAlJatF829QBtaCXfnbH3WV6Y2gaPiHVY4lQcv5
EPt1ZxXeteQ6/5DY/WhY5IJGouncb/A4b21z772Y+etE4v8oaGDJelKX75bFWRb2
NEC8uh6DteOwZEPCAy/2bngAjxmZvC+1+xxeXMQE9UeDOZNGkdrVHKS2HZvDMwct
FhuLjER+vMHr37I6qGMNyc5uOC2hdsDRNuMMGBmHXi6N3Q5yr4S1iMrwKe6ZcKy5
6jhrrVVk1w8TcjTUslgqGZV1OlIAS3GEMTGNXghZcAUh6yluVRDoT5DFR5tE5/JT
337mzaXrhckw7lsPcAtWcY46NEg5FgW058UmC/FmavVYA9xOjJzxYoiga5IS3Mls
WqNqm+OaxLiF4ldH9z8xIayDmjS+c9andVTE0M8mDjjfeSVnz6tdTP+r/Icr5W4u
HVt2MJLzPZ0Cyk4qMCB74/wXcStxNK+cdQp1xxr5h4ZfwwmMRsoLtj4Gmx0dw50Z
EnFwVYpENsk62q+JrdPpFExEf5L5f16430R4aSkvdufsbfgnv4tfjNDOA91i3eNx
qPiq7S6HPIGBrG7zgPqmyE+2SYqaIq0Ab/DcH5WjW74NJUIcjwRqvLa/5CVqIxPs
4GDV14O71ksBZfPybIxNgiAHK+3Ye0rkwuES6eR2LNxJeBINrwc+nMI2z9ISumzU
5EzzCdqKwY+ihp1uRfCmJLjQ3Q7HGZPd5vBiUXgk5gLW6R+CwoGFnRRSLJmP0Pzt
PXqBjT9CxmMt3I1ZAhQMmhvdPkDudLZPwf2rAogryKE0FRciUTsul7AilTTEcNgA
ngFUSqrPcEOqY0x137STykqTtSlZIftnBd3Fh3poCFf9Xfo/bSA5DgE7Y6g2KfNc
4UTinA+JywyKFoxyTZWqVxA6DJ04aQX2PWl8w+kaNgh+pxjcmgSExZqb245qGHDB
MBlXP0RMTdi4HEsALXWBy04ZH8YlL5Di19bkxIIh+JEhAxbTQtl7UYZZqx+yXA6c
w7cyvu8rE9NHS21pJBAdYwTPZh0giajfwrjqjXeawdOdBbqWoS3Dy91FyIre4NLB
BKIoLg+Lem0Lip9o8hWm20y+lejYJsSUETEhL5b2gPIL8HMaJwJP3P1nJHj8qNoN
Aag75EpoXRK38n0EiKoElC7Xwe2SIVmzpl0N4FQQWdhy4uYNuRalhMjxYLPPsIqX
ChvGAPXl7OeawbKgSDTVfqXXkjuPrgJzRl+7whi6Eng83sruzsGNV2hjtpr1U7mv
tNylqbrrbkVuT3qXLPD0AAdz1OacPw+82vNOw1mTz27FeJjRmN8DMTWI456zv576
iGL9iEqfl+VxF8f4HCcEa60OwXWwOc0r1cRCD97kQyx27NV0SzvWhTzaJOK+xZel
OheDT4XpquiGydLE7YJ/M1vU7QSkH8m3Orft/PbUJq4nlSy3Ohu4VisxWsrgQARE
WO2f/KKGZhI3KYq6PDyVlQT4ICCjyX7H6VO8K9C8eDGJpcEoxa8eUzKiw7WQH5mJ
pbV3GC29YEzNjl7bVi4lCxe3GuRuuNFwYrsFewvZDyx4CxDG2hW+FtkGCYXRqrlL
qqiwDOlLpBdyWY806LwC7anaENGtWmesbPbYOevJ9wdOBO/MjhRnC7m//dkCNw3S
tlN28FMzrSQadFVhxcLWiVN9motfJEKpxV0Xv+Uy/O0SmANw36SSDzY9fdivREYw
o9dRGPk1SyvHlMMD5QOeoh1l4WFq5kdpkYcyAyamAzhOKa0bDUhKDHipqecgvcBu
bEjYL9XSenkOmaoHS61rzjaJx7jRgdQRayZrhcaN5abseDh3AEN72cRzSedMgDv9
5wPGmvXYnyHaqn2PdaHi3zqw/EwSd/SpFQrMcBGOM8dLfMFtDNt4VBQ3Qnn++riz
IY6fulW/NDAHDs5bL1cZerFYY1BaLkNlQLGCQe1KHqc8x+dM90LtcVIbLzjXjFo9
sPywA4swd0dGYuNQeNuNhbMVD20mSU/qZ2Mwfl8uKoRyiLQHm6e50KSvxB/ZtVp9
W8c7dQOljsIV+kkWaxPaTpaOQ37B+S8+Kzm7skUSuq5qu1q8YW33e/Y8tGiegW8Z
pZ97PEFz2pBOZTtnGxSGObqPKpIRMkbk9FpqUaGIEf+16WCalPEqeWa99EEBq7UG
ZPWssGczKI7CK7k0baNEVgKzyMd37TcrlJEOKhGm8Q5Oze8Qm85KsZjzXAUFR9sA
8+pJByZERtSYFTA5dZ0C1k3VQ4U+J32Rop07j6PB5DamwjhHSzvpf+k8j0fxXqtC
5ZCWp9uCIwhJHBu132tpuatiIhffz9VvuMrne2uqd986DIEssG4YmQJ9sDfv+Mr6
OFTCuwwhgcgKaC1nU8UuwFCG2jlnBMzSFloJ3MFxCnwrxaVmeECyR1yRowicmKdy
+9C0MqGV74WTakx/BZWY/0d1pdhj5kYEtn66sLFquhGFzXVRkFBqCsmHL07G0oxq
e+AYkL1TphfjsZTjJWohCNswoWi4WOd13vjhS9Sw4asMlfCv1k0OPt1ipO9gs2Pj
2j7l4J2yGkGZAS+t/UCIjEYYNETMIq3L+qgYDm9awDy3Z5XbZ4ZyadYVdtXGCQE0
522/PqomXw9hr6sCa3U+X8mQelCN05kasiMz/gNnjySBO67fo+kG5IaWLy5eFThV
rgM++9erlbS2i2++c7QNbvtoKEAV5J4kP+b5tLkPgDYVFtLzyLuljm/OsSdokb/0
wiwUQlYB9ZBQD/UZeW2c+Lyz9uLlsJ3WAbQEPDRT3IDq0sWSvyfbO0TQkYN3rVAP
BYTldNVzSGPjjqG0Qq3EOTIXeGohLdUjjmDeOrHwFP6/z6WpbrkN7dVxTMIBpe6j
DSA+qM7oT77vEiM4CB1To/e0AmhgnqD8Y9AnZk4wWy1quuaGL26t2p5cGfgcLHGw
ufBcRBYQf+K/yPSlDScwUF4yu3FFpvaJeqxXh+ckPjum6MJUiHjAnKTJbnBJv3/m
Lk0YXR6P2KpeJqx7ZsuobLmQzt5fBCsxiD65gq4Kb8K8XNr/Fm7cUnfCZOmyX+M9
ar8+wOjcdizyz6CImtYMSkgYprvTyeEgyLoa6h0U4JBaSnWkg4B7u0TGYYLJS+3I
a5kmcQ8ViEUgRFzM0Xxf5XCevuWkn2hA6l9hq7woQg+i2PbWfI2BBC7UKnXYkA4v
VACY7FMuH4g5uFIJq317ltMGKPJ0qdOt5j0EHjkZT2wYlKjFBU5IZgeC/8UfEZYZ
LiajEreFo9J9K6a812s6P+n+Wku2bQJm2uw0r5hHwg4kgZo5+PqET+CV5jWF57tl
LwS+RNHNDvMMialOC/BD9iRX95twUUty6jq/eit7M2hLFVVMVkbiujqvIrFsya1u
aDomH5pdoU4FLcAjLIpJjS31VIdTWASIc5U5HraXQOThbFyMi6kB2ECibGWC2NoW
MElZ0+r79D93uQrZ5VSuZDrWBfbVAY8M5u5N6NIABFSBO2rchoSvEbYZ4m/E+8bB
tgCSRDwZ5jEEDBxl9KeWyUuC8paoyeaegrxgXiwPOGmOwfRdUQG67a1kIYVr+ecN
tOtl/uEKbPdQxNaGswpyt6atik52OkzArrVU9RFol4h8rmvA74i9RVrX86rgzF2N
3NxY+3sGYiL0SyfTT8gA9Y/zKpuVEoOzjJkJtlHAvRggF1U/p/qfFML+PJZwvhq6
OTtyBkUC58OtIGmi43/Evw7BFeEWfbz+a4R3pVp5BVNzF2FYOF5e++C6Ug/3D5RY
16Hv5jh/zfOeegVk9usJcAxCwcEFs9dmJkn3QdRSicnS5F1X9p00D/1isdMkp3h2
Wc7ISVdJmEWpgfWfJydeSWkct13r7a+8LlRxrqxcvWQMC+ueeLLWsGBC4S05ZcKD
dJ+f2L+64v8mZlQUIhWtMop8lls3YsmBgkbhKKQU0r7VKD6zQLMTcq9Dmq/wUJM+
/06DaSRajB8awuHe82WVzr202Xp75X9H6Xxw/R/0lo3tiq/FEu3mjvmH+kiTI1/s
uxhLhRLsnjwz4V8GswtZ4sDlGSCLiyNJ2hiSF3f+6zLL6CXzTBIQnQ/EtrLqKUs/
ckNZwqAo6MSxAjwbX4NxbP5Kgk2Ns8kE0M2Ztq782Ur+iFMmzzJRGTrX4VG2rG8m
R3BOmbpz3W8jZeXLEO/BR+AX0oEqwBxI5XcH8lnfVORBkOU6iivVgIh11AhA6A/F
CoVPSjU5d+8fwlEzHfV4FMH6nvJzP9to6v+7DspkTLzFQROMeC53PVRgMDopcJTz
NFdPavu+AxARoX+Fq2a7P/BgO0CSkSEQSMpFRpDb9DqPaJ0rWnRzPO7YjuunbwxM
RgTSKkgygz9dDj/3JUBZqbvr3v/tEWl4kqCoUjX2VPD4uR7dEgEwuNcxWT8SsTmU
YIkE8cC1u/Kfu7+XReczxZVWahaORl+wZ92oLH8Ek3C+DGm1C0/f93UXuwN2SXHd
/SILFBWccwryQzMi6NOSs39UBjvSYBuaJxvW2ePA5jPSq7mMSfjdaXzku1QsB2Qo
qQYx8/3gU6CmzuAXPqGGvj4fiNqWHNuh2bRRti2fx8r5SJ1fltZRWtkap8GJBnOl
FUZpJ9rxMpVGJjYNdxtAFrbkmFH4o7hlrzisrCmnqQAFN2ZNnGJQpoFN0Hsxh7ts
uUK4vzdFGcValgV1GQz9MEbimVBRl8DlvDGJ8iTc5nJERBOebR05fF+pAT+2Nb3l
4XrApFSOdf7vh2eM6GhBeS2uhLYzunPlCXMqf4RJN9fLZChBG80CxhxTdb7oMxPk
+KBF5gY14Cfzjca9Xw74rIODm5V6VZO3jmAcO/1puLnylOkGnmhnUwV+Tl4kLtya
IW/YyVc3wvXkMYdgpK88tTm9HDg9hNJfJKXODzs12FEm19Lf8xB540ZS7/OEm5zx
PzLehE82jGlRZuyjif/sEwZuN72osZRhYuVe+VwRJsg7lXD3SFV9lIhoN++Wuexs
dAwEM2SHOatIvjyf7GKBXg4s3yZe3qZP9eZP5YuX5yiwrHLlC3IPonDYc0yk8FPd
Q/xcYB1ti+lSrPW3VByh9ym1phSsNoSZcdMlr61hkyD2ARUWZwoJPgxhbJKaa4Jv
ANRorDSfoRcPXDdDmkn8C8GO1ATvfMInOhK+FtKV450AlYTY9GcZy7y0pU3kS4jd
bElkg7MXrM58rfXBDRXYUpbtrcnATnRtK5Emdx3Ezi1mEz9t2mmzr8EPXYn+xxOc
o8eUzSm9qu8QVaY/tHJlxyt6ZmRY3x76YJNBouSpoS4n94LZePwwHH51tHTmNvZD
vG2ZDs6UHXC0tWuToD8hWuBMIv57Q1IkFBYqdHuVTbLn2DD2Un+uPwk6X6H3A/O8
HuSNmRQaE8frQ751Q4K2nx9VrDV46Wx63n6x2DcQ5zeV7iEkoHQ7Na4utBkBBAJP
zwAw1k3VrXicb/aEWVllV8fe0cocG+f6OnleCAL+vk9O7LATf9nX+isIj8iP/8Mi
byJXPVKaz+wCrLP2qsLNZBDqOc2PlsSp3XIlPNDVGybJpAscMEcguN2L31mnMzx3
1XDNs0gw1iaF+66Ai4YlzfifdaBV8k7ExO60/e5WYbZoJjJVrWcQcb5mvfnf/SO4
3r9hh34OqxNgvzxWGUWrrqnZx21OJcc2QJvtwkc1A7QLBv9W1YBNR1SQl0sBK1Mr
fnaRN1BxuVr7pNY0GYAmVNj9DcUZ4yw65AdVuG6D76x5+XcP7FncRBdcDrdzrbJS
4bGYRZ/eVP7Ul/Mi3NB+NuUM2PNYq3Ykrvb/Qt2bXNLAfqwKg1PNk6ZIhD7MIGCS
6F46qMaqJJEOKRCQE0alh92Wvf5GmBpovcW8QtEDypdvXhU+cfxexGikaqWIZ0/i
qTSVBKPWS8UttZ3kiBemowpjXXuPDGVASLxQO1lKFk8+XjbraX583Wi5rXfHsrl+
yCYzkH6rWHMKFlhJlz9HADgw8gcSq+GMz7C3KDb2aGzf2V7B/jp0q6q9guivsvJ9
alhFBsjUXsDFS9Eon+SMRBvk+xa1DkjnLGQROYIYo2pm4cWEYGbL2yv8mCbskR6M
bnClLn2zF+9NrDJyxADF+EvXJ1+Xi6BjkUTbuPGvQw40o2pKbvZMNj3CPDzI+CEf
lDyUVzjT058JdfLf5aRnRhzglQ56tGD7LqLYvzdX/jb7wrMwclQTDx24uh3oWeBE
H86m+K0iJn/s4scZPs3FO9gFkibCRKgrWhaYdlShCBeHxcoeetU45UOLOs698xow
5SVgSzT/u1B+mCtbEHLeXlWBf/OY2vLH1lr6DFuTalzd609II/4QjCEI41vYMEfb
xHKcUlxnq6F5DK07b4//MxYn53Vq96GpRVAAW5NoY6EO7cf9qQdPwPqABDti23ZM
DqikPLZj52TnZkTRiW9IqgBQ0TPd+xcCbLWFliR7gw4AsCWwZWvDT4oDC/zh9hr5
AgCTRdF31WijlYJ9ZHSAcrHehBCOeu7A/fwBPVYzkarVYYj/q1qsx7FDcWaFt+X9
A4p8jHKZMSpKVbd/Eaz+JXjZN1cselPQr5STGrBjFaEJ/kgh8/otY7Gh4jL6dT/h
XI+Q45CIVUrkLAiuHt/Dz8HSpd4PcuG/PTG3iG5L/koO+tNfCD+AixgsxUeNEGQN
hS6ASjxwifxgjUaatOwnBu8L/YUUaPI04I3LrubpR3C9puJShSk0SQNXi9Cih5vQ
7td7gtWIADhgi+DxMqnEf8IiFnhWfz2w2RhS0SmIeN35wqktVHDkVBHmj70WQ/SA
wj9EMOw9ZVqhR6sYtuCBE+nObqYPhUVLAOrBpX3PlJDbUUAqoxtGf0eGdz6P3i4+
t35t0cuVUAaKOQVnhtKppNyAP0isRHfjbvlxmDRb+LYAYsHHsrLAhJYW+yUKwKPF
3B9qsZHB7lzZm+m/9ghlWkdlauSep5gEZE8SNH461OEIORVq14/9KTs57XqMcq61
rZuK/O77Dh+XMVE7zoUwRG8I8VFoq/H2rR63VUqUR3NdqAkiuWXBN9MjDKcMUhsi
ShQbxuNj9EkBUNrY1Z3rDCqP9wgoqNtqzVcAQI0Wt69zgyHiJ7dCDDHlIoLA5bhq
Lozcd7cv+dBL0XYIDPJRIAosDCBO+RLnT2ldxIRIQsYXf+KrvT3+nsCvPBcChkZL
zs+6ewfyoYDj15u3qbFDI3iEmxDgqr8DvFFMjPPdRAyLrwrPP/B6zmU8lzAgL6mh
lQHDAgVh9oG8m3CXYnbO7JnV1LOJ8p4DeIknVkBrpuwU0uOt8exCO5O9k4TqbZGp
OJCb753UUsuC4NCx8QEw4O71ZsNLxdasOsgPim1S1r/7jKIVSiD70w/zOpeC2Z8H
yBLYmCb85Sb17/uGNNm8Qhj8a5EVx61+hMf3cc5Wq2xtfKRwJkqMfvBmd24ddLMb
iZGiio+jsh+ixr/pVEHX0TK3iqS2LkWBbzTEvbtpa252fzL4wYVNKHDCd9elFAov
kYXnoorfGvU5sfO1QpFLd02bxGlsscMXgUmcqg0QvV2GRiS1LveS/AUoLLi6o4cq
kNKUn0PHx1QpHlXyoRfP5ggdPfP6eiqf9KLKjIhs4smewa2EO4KihOARyn9FNZBP
pdiALxuj9Rnj+oZZsYCBh5G982QhbdszCXQEA9Nr4+vo8IZ+4eK5og0HD2+SIGDH
62vLKcgur+vYJlb0jRNUjufnUCBo1H7cZlZRNLS2V9RzYtaFsgYE4Odik91rewHz
ZdD0S1fqqqlMHNhCz9eOG3x4xO/JX6jZsm/+7eFXUmqK4a/W0ApObxjy2+u6RuV+
WhzZdRvvPdoIxjmkc83gp65jYJ+tESjny9CojY6lE1nmf7lsaJjZbSkndzptFobm
/j/bACSVfZYTMEtpos7hKBljLGy2KcozJNkBOWt7Md/6K2r4dtlEc1IlALjGwm2z
nCuCJpQ2tH3Sn49I7k2KRmWWCe/XN2RuqhsA0ZvsolvGJzxzRcClRbYYfbgndeEG
CWFkTnSPSv8cG2aBHbva4da2rdB8wH/WXrC08ayEMzhPcEzXabrlu6hj8zvH06kz
onlwE0ZkusvJ0IaNRyfMGJnmpc1hrHOxCT9HdkHCiq3A39ZE4V+KQgurF1AbuBzy
PDZEl6vRdRbYSPMsSrJy8sjmWePt8J0kx0vqcoBJF2ZovQs+L3RyxbKxEBXrYSRr
k8ahEzPxuyGygKpEeS21ocsgA0cmrqXS9oYuE6FXRyJmqWpJn8EP1P3ohwyN19kh
zkLdHXOMCjq7IuRCkkBccEqa1++fe9C0ep38gsrTrFBhvJpjVptyRzyyI7Ds/dLx
1E4xVh4nFhXHMGKuyeBQza7aGLh2hMJ/M3muXuKjTzYB1yzf8AmKPYRVE0RgeaYu
1WTNukgfRpBSnS5jEli8uLge4ZnTtFXr5wmUDToikatCmilWxpz6358ZQiEQ1NQV
1xij3lXfwR+PMnDIpd8PNSInrRspY1Lm7tOaYpcvO5XBhV9yEk/yPpVzCFEpIQkh
rOm9vhmgPiYxPSflZinYqh94lmWAteISVIQkeXczeiQZzpUt4T3WpgXBqNdSWf34
nX5WdxFGLEKax3rFJU4mW03GS6LrqpXqQ3rYV/JJDJviY2t+KS0KEvOirMqz26rX
pg10W9hkGYGohti493h4/g/AeLjGi2UfDqVXAxP19sJkzqnY8gKbE385up33tACI
0qwGYe/0K+n344w0wzi56OWCKUR0v3Fvr4QQxbbRYxXSmpwsYWOukQhHCqGXssWg
Z/fXf+qtTKPwpyXfMsbNMnVvgELe7t+hoVSkm//zBMFSbW8303Z29hgAnRStvUUJ
qxNb7B8M79//1aVysHGIwCrnkLGviCm1hdnMH7JGNIK9Sfa8+0/v1/blvppWjFM1
28t6qpud8AVRXMHd0xYBfhsGXUBMEQN4q1guH6Cfd0vsRjRepJ9vvJ9m8Rh2HcJz
LenGhyj/5GQF9MgZBLM1d7GwYOlUEEYXdVCI8+lTeVI77O/5TQaYUmkmQoANVTOg
JNtMKStZJ0Xb7OCMpg33zcxV5BVMJXTY+qb8+i5PpGctGmVXk5QR9Vxv5RyQxZxG
7JAyMFCZ8c3onG5GvzMUq6sR/vrLFEO1SoE//7j82GK8I+/oJAaMLVMICISRe3Lu
/Dj2oTOp6yZ6/3mOJNa3fWb7prr5QpDBdQll/IBFrpegcJxkJigB4l7KlmSRFRll
5/5eba+lq816GG9MG2NhcbwCF1yF0xl5Xq7jdTQP44mzL8wXfkLeAl36BIJkr4RK
72XMPgsi1bpJl5mTGVRxL/KdHS+cDI3pymODm9u+q1jthd163/9xkDo8LjIVGUig
RSgE6r1aMzjwCfPSrjz9rBT1OCZ6JSpTyHg6cjWESvFP9pTebT2VNsmqyrUOpVyS
Owp4Wha9mAdli/o2lYyeyw5U+MoVAw+sqSrsi3sAqaBLM+MxtEqJnx8+uMuALKsl
+6bgqonN9+6AVwuxoi61WUAW4MvM5HqtN2J0U/lXY5qkF3btFSOveEfhhv6RHkrM
ySXSIMt0TSmPEUnpafGtkG8sFfV2oltgs4SgzC0uqfwNZMdnGCE932LJrNlMVEJ+
WyTVBpzjHiwpO8tXsS8jhBUsvZemc2IjmRyydLz+EOxjnNVA8PKsB5tixYnspluD
qU5GPjLX0v9O/a53F9uwSINKJg9jSmySWn35LfD0MzPl0VtWTnFqBd2oRiid/9QV
U6T2jzvxwJGFseHlFgzvLsdhToTzox8GK6qowgBV/Mv4tRLyds0r8Ic0AWjMqaKq
GhOWAbE/i+5smTWgV4+WtSV8QO/JTky84jqJ0UdgoZSypsriHfvFV98ZiLmtO3DD
Rv8dCYlrpmlmzPXJ7l+fbxLPI+z0PyNIlnyPZvH47VDWKsHv/tpiMee57iOTqU9M
arOuQgNdb473bsErwoPd+odaU9ySwowFnmSx0F8rXp0ya9dGtSDXgJ3y91zSLspI
XVDOv9rVGqNkaWhowrXF3jQ+mX8M9j3vnx5wkgrK1SxIgF7tEu6NYi7Y+I0KPm2J
e4ly01YxWUGAuIkeKwYMuvD0WsVyp2psEagP5iveQ5IKMWin6rnjRurm9dQpOmD0
W38gtadF0JcU/6C2j0/T4RGkaY80TxxjqM2TJv0nqagIKXki/4MunfNQ6llvcLUe
vasxMXR8ALb+Sx043etpO3rW+h++chDvqkB30V7w02IijA2RVQKTzXQEnwv0Ru/h
Fu4jh1SFVBaQi8qif7HDt8X6YudmIp1xD+mrw5omm1Bue260RiKR2Dme70PljjpF
wGlsB+wD6djSJH0nnPD363KPfRwKYh8SobdypM1KoUNiyPK3q7UDzcW2orJ/+a2p
MdjGqFWbIqJKipY/2RaHWYntQl88Y27+7RqskuEdhA2Tk0v7v78R2/3OxBVSSJj6
njuA0TT9FB61rnkDRiuqW5Q2QSsTAAMiAR4y4vnhgTqAg/fLeVhYo1AsebfQbJhk
Sk1RFBFUexr7tz3IhU2e5gLdNNxEqz98Qys8EjXMnZJmzdLlOhk3haXB8d55O7la
1yR4uEbE5rpqmPx/wkvuLm0+UZ/iIvwyb/7vWLHjEY5WlNw107fGeaOb4tW8vcYq
D4zXKyFCr1b3b1dmmTN8JjLeRnhP/fMI2MKfxvkg+wfUg9Im11EDifAoMXelsfI1
q73BzRWMNlsnSO/nFLjzJR7353SZFwrHXZ6tiPR0UiVc/zN0j7JI/o6LtctdDSsw
spgApMt41pLfPBOt/3jpk2PWl37DGQC3YCl7DrBI55DoL9g4RvjU/3H5RhWD/Pqe
L97PgSvMwdQwjku1jSmKCapJiAJmZvCyKTeuZBGYMsfIXrAyoxTzyrGU7bd2qgE3
LQ1v+3aZQw4oVxVJCjiJwoRVte+PhFfIaLqPsEQy7zUsonS4IgYL5mQRLsxac8ml
Z+n2tvT9rPIxV4Ha9VY9PxTNLQIu+h3PGJDbFSf/hY5XzB1Ya/2HTVS0EKNIYuDv
R94TYmZmJCAM5vnFLDUufCpnwcPfdKYQl2Irq4FKcaT9g1Wx5gQA95WhC3Xm519c
sdXK36V9/U1FLC/gVlYJ5SrVxovx3CCLnYeRxarJMekSFvvLEWwRGTsTWCbSDUul
OpLYuJwBWP/J+Zj+biYG6CEyGTwB86Y8bBlSEUrLS6UDUh2vzQuXILcobe7KQXgj
U8sPaLm/W9LaWX6vSfro6D7EbHOjAzfT3bU7I4IkW3PDmcEZndQ4gMi12hUITRmp
/PA0pPpLGyFDlU59bS1dNAEuo+8VhV0ct30W0qRLovtRge6zRveUCTamBN8znwFr
NbAieIg7v3lj72ePqdv40WO0jLuvIR5IAndRD17PbIq5cNjGF2PFEQT00Id2yNxj
S1uwFGsT61KrczL8evDQEpjDyHDhgf69EqY7vjiOOtiMwNR+SywCmjxOL7C4uUB0
y4a8eFaUZFLs5x8VlyCqEvc6xiQ4CM6eaEfVRiLWldK8kZ3Hb8dQCGSy54eT5UQo
dL9l3xKls61LK9ksW4m2H/XllxaukcTv02sUDX6UEYXCH0RUPg0j4Y4N9wyCiEq9
a8bCQrfJfVQP+5R+us2lcs8Tf3pWw1m7KuEnPjkvmly++3tyAWN0X3hciAt/YGgW
9c9pf8kXtP2qOs8mGXjiEwlDrlsZ2SM7UEHj0pS5RDVim8ldxREWG838hLuYnjAJ
j4XRRG7iCyNR3tH0ZDmk7f2CxnIzU0I+KnmeURkRBLX+hgFLskTUelYh8SxXsZUT
3zdIgBfJCw9fTsVn9G8QusJR4UQInkIAti74EIdZDVKtPzMtgntIPg3pJs4EjiiE
n6I0sMwbA6maYLRdrTEwj4YidwAcBHq2u4njp1i3W5zGy0PNn5IXlP1QlGxBQMch
I6gxE/FMexBQsT6s2EJ6AevJ8MEYh3pzfY6dSxDc8aHRupuAW9s76q85tHmu0V/q
gL9O9/gxC0rcxqdHijAzcLFSW45jCrsGGNnHm7WQzZE9o5bDr7K1RK4aifYvC5wd
favCJAGqKsosH7b85b3cKytdajByKoAd11UYHbseaXAilpqkLN4e7tXrmO+d21+a
HHEfpn+D2MAGQjpbvu0TDjfzbys2L/bnSuCinSFgoTKqzzBfzZNPFJsmLK1mLeeP
og/J+ehG0ZZ9RIXFIW87pwYcYA5W0KK3tKtWJkf1w9Um/0DyqeCCkOnnz4ATaMz9
UUkRNfiye45wkOFAKcUFexnPSvfvmk3cbUCwr+7Gwo808gB6xlz7iUdMBlfacv+P
hsqGDqn+R/PpolPwsRufqclSquIBlwrc/06Gxg5hQNiQk2IMR9xlIM5z3CZX0ga4
F3YLAyS5b2d+eQlYk1xQCIDDp6DIu0mjTOuD1AlZS60BDkpRSBvIb2paTuHANfe3
j1+Ixd8cyXxI4LskGFpgj51TMnP0OvzgCW+XSRZXFtA0BNufAeJNdM0VWg/RIyJw
zRhjynjaBrxYv+wLyTReUWf2C+xRLdr89oKvKYCOsUmKMvM4wepDEGjJckdTqf2X
Iql8723OUx2kluhcUngeKa+mdtP5iNR5/k7MkkarxvXiMijAwjC7fradePAunRoH
+CzWfO8Iome2lPBBlfvZ7SJoLgd/stRy57CsC3IdifzmGb9rfOBzCCktqgpUIgKE
enbdlYn1EKbSomHaXEJPpoj98UJFDuxEeoEcOF2TxUfTf+kk4oEAlhZJxodaG+zI
r1vHI5BJRzqkJRUW4ARUAZ1+eJ0lFkFPi5OuDoppmWQpIkqWbiXJt7un1rTCs0bl
/yaDmm4iHW2OkWXOp7YuF/Y/DCkHZIxoHg4KESg3oEXTuEd4lLtfiHq+8RDXLHL/
d5mUhe+YLFUxmChE+KBwEMhBR1zusl7vyRr/FIjBDC7i1CYLBnJeCVsJhQX+jMBz
wOim/38hUb7cLJbPg5czaV/cSzgd4dKHHWNR8DcCKcDYbHhl4cPVWPcNCKLz3O7z
p8jx1EEeNGpejTMF2vTIIZGp6sem3DbgXLXSMmcks7G5Iv9ZJ8VbOALp/1yJum5r
dpDynT1DNGI+Lk87QFVICUWhMvugtKdGbeEkNUxv33/3H6STSulF07OBtVlg3IY4
pAHriCxjriHPqWjth5kGkZqzL3Oe6jjn7gmMrIZEBHwCZOagVAjBh9QqatanrG9h
MRUUmbkrxmyMwF5U+N+BXK052NRtj9m757YEnaIggY7JhTdXCvHDsuLr1yjKBVwi
qdtjiPMBvg2zmRv227q7xv1MWDwECYVcQRyNSkgySnm0Bke5F93kKDSKE+k5jwjM
kn/yfN8+iGXx8mV+4YrOMn0DuVLIledPSBYttqPtmzN7YuZckWo0+pTCGMWSSTzS
c1xrPFNxSshk0pXUkhyYJrY3jp72/DASg5x6jPnm7Dat9KvfPEksn6/a4LgU3w5f
q9t/DV3RIGLYf3ruiT61+pO/UT1Z+J1VwPkshj1YRUJpi1YjIO440BSdRyY2CoUz
D37WZWzV0bubdakNDWM/0rGIs7vMauv/1wvOXQauQjlnXg65zb3vlnMgyRWIIdi/
tLoddAe4tTdsvYZ3wNaFH+pqvp8xhFpbRVVISQGfoRkV6MnFguz79oYMdEfb9emh
9eMiJm7DAQfuyRyKx1kJ1QGnMyoXPpXTEez5+CL2vtbWH+9EZz61l4NmPTkjCaeB
YXEKVbOyizpN4PjzrvD9KKrE5cHA2V17BrjcZ54R1iIOCYCHjAVceujYk7tOLflQ
q8x0kGpEXLOzxJWCzKBtnxOW0pSnYuTd6yv7nHhcmuuBhwBdmqj9gJYIpdDdyb4U
rXfT2tOW4bbPiNNR0BN56kOisnOJM9nFJq+HWXoQtYXSGfem9wayk9o6dTZE9f67
JS3Lw/06NhfaBewm+wsOQLdQkQobpU5nlBdGhee5yzuB16tXK9iS9PPrrTc+sT85
KlWf6DGdF7FG3/ViJN3GO2xtfML/MLZQ6AfjR5Y9nltuGUD8404OCnyq1/602F3t
uDeX9RzpEbbslJLbx7eMsO9JQX0hITx2XDBCyMno0GqYyl8Ar8NYZh4uhB0cL2fx
+K9jHtSVOXZc/a2979eWVYjqScHAAAAonjnNk83yMjHx/3BnTK83bNPhHFdO9ZMu
nW0+hLjnb5axGeTfdSjTKvOp1cBChu3u7APl67ghOUa4mutqBrUAN6/UHrfUGMT2
hjeM6atPLeGPNj5nrIu4O/i21XJjYreQBBfeKNXIW0gu773219P2JSFo+03qrsXC
38LRYoyuo8R4XuADQZJR93pUnPVtqJ9qOV8hnnuVjQlV1mN4TyykYlGjpJ7R9mk7
fo7l+9IDX5Gzx2fj6qZosBveOeLa7Tee9WfS6fLlIIuVErgPWpw1+gKVxkw3cnRn
UtoIxGws6WJTP5JNBljIhseUqaIf0ieW3sP7I3OFE7M7k0nNDfnhC3HnufcB35rp
l5BGJdYLnuAHjp6w8WgB2sNYn67IOdXvNOy7pVNB52HD1P6eRUve4HLim3X/2Baj
FZEUTY3SFP3i2NluCFbCthXNXCMBTvj9Xj///1Gp4YCHQv2f/iFVPilTh+tFDYL2
+XIOIrx59S3UEmeHlPrQlV3gALjsG0RVCYwPY+nLUmCoVqhH1u7SNPslTGc5h4aY
0HqJAbWfv6V+hfwwSg88Ncj9zKRcmbd9alVpR+2YQ9glKXpD0954aI9tmoz9bDAG
szSDJpySgJ/3LPRliol7xQ6r/UAFwYXpF2E/izz9gsrWbFgFA8tCPkvb/G8gAswa
3fkEox0REDi1grTmGoFXmg/68i2s5TZ8IPqxmAF0J+QPs1+8QwiQOhhpAWVKt6nA
olqYDj+k9luRw/K5te6ltEjVPRfNs3xL+GSX8ijan+mg6+UBNNVMhMl+RTbh6gDu
ebC5dl3w9Z9LTTchT3+WpOVNsCymdCO9bLTLjUAgwhP8Morn48GveIpYWcjlOys3
QBmMlMAzfp5ErA/gABK//q4f/kUL4Ycco95UYbw+nMJ3uvAsnlHtP/4tkWC0XRqz
k85ZuUGPf3SwURczCBHCuv9jPhEDLvBCLWT2tslGyM26Af7mlQF7/rz0d3aJ3taS
OTeQUyEpVywkBzmMPOsps4M/T4BzrNs3opa5itapYE16sE0TCAJhCGyM8Lac6smR
fv4ptYstU3Qxbn7YVNlgcQobe46p6rtZiFrZ8cxOEZwBfuSpisLDO+8QD+640xR2
+THtFFtLXD3oPQRWTlCtGlWjz7KHLdbeynVHl/+QyxnFDk4XKYAzZnw6A7c923UL
Jha23pQk9XrW05TsrJ2uT5tJ+5ZTyPNJ1dwqwMNSMR/fTyrNgn4a+yJTChoEle+q
Nexcf+8a6dI2tMG8B6uaJfJI7zDJ3PuXDzZ91NYvk07KOu08d5W3fgz2HQaSFqYK
Sqf0tQmq0YOhEQv3OUytfsUUM/4PlJLEGVfxYM+E6luhy+Ht3iDLoV2JW1w8T1Np
tw45qNUxoDG01Lz65BTe9Ua5TVd8kaJ7Q8kee9MZryepZ0Dy0YAjebGiJaJqQ9IT
6uIfrWGHDjp1F14VYp3bHoz7c53lvpMWXFvivyat4Qdd5Rj76zj9dpwA2sqjIXCf
oZB8RYY5xeiLwOgvwmnIYizyoUII/tIBy8UlEikJaywI9AzoWrxs+srF6s/o0PhA
MX6JXwLrtpk5P7Zt8CMqE/6vKLloOnRud/4sbpVlRv0hYUB/EyzLhint8e5mcAS5
SMyBimL3POe/mN6ems9i0DOwLY7gNvdotyOjHA4/35aQmpRY60thG7u7EqqqEGj/
9axfFB11Orzb3T5Zmfl/8V0gT/ZYZsxA31BZEGZJH0QGNSHd+grOAtmNMsRFxTnU
Y5xHkpe4M07s2Bk+XJkKhbGkYy0/XmOqL9GIily0BXVxHubFBgKg2Wzv+CoteJxY
dmUfdabTQn144g7DIP/gGJ+aklZyS2ICuvm7xM+glhKIpSSU6sDbvdj+QsvqF15h
mffJGtnHm2gA3IRVOXDJlK+7mbNMxTP31BZXRVwxPrNe4cMTaO/318n4YMfh/3B4
fOd8rRUakJtiJTzHpYT0wskv7lYsdmVXCDTX7BVPGbpRYUYIMlG4bJtLsacG1rg2
1RzsE40t2nyut2rh05/pR91Jf5DTVvbb7e+4yebvt+3iFocVVjmFLrFHoo+Asw1M
WPJHal1gMtl42sMPnFQJA4QR4TArUBSmScLVe7LTTefyKW2TEPiuvY9IsF1R8773
jUYoPXfqjbVuyt3/2mVKBIu3KYZjsiUvc6FeCW/q3uJ2e3noxysOJ7hUWBbut52J
6VrbVW1zMMDwqIlnVqa4W8pJ+hXf57ZS24QPY4+Zm6Ii2LIZuhHwCc3FbGpTt2s0
E7BawOdjdS5MKNxfcBkcQ+sGJhP/XKqgMLJC84l8QWAObtOx3nSXGP33Fmxo+Z8p
KciSd0cuqr23B3tw/R9rTys8QjhEPHAuz41gcxDJ31Mu/5mhMPTNJAwwSQ2QBGsb
XJ/uetzzesK+zQRR3p52hCDA+nA/mHSQs9zwD/HoNK4/IzwS7OZs4Mkxd8Q1tN/L
OuVf1QAb8RkCY83zGBZ6JARqbje4B4XqrKHIzWegMPv9S0ltNEx47lD22V/OscFC
dWWCADChMdX3mHSAtdahMXvO3GuoKMjXH07hEuHjFMvtpvSN2YkOZ4ZpldbItWmD
9bdxiAl04OrVmxVHKu6G8dFQ+tfmMJ/+GCKWRwDhq3jzHiWLX4D9pag2Sz/1qJe2
CLrFHuVQiXcuBRZKgfR0GA8T00CZJJUrHRyzfLzUWK/THn0raiGiqDkzKiLlqGx3
wrdN7X8lQAAavvvnUIOm9bG3WpiYKQ3JrT3uv+hGmjDKyDtF4faJWtgg5dpsSwAU
YhNPnTkMGryMY4LZ2vUgon481ausESXYXEH3k4kEol1IfacJdBPWOSSbnzHls86u
pWKZUOc7Do16VXX1rsZeUhF6uOalZJFGDvuI1FH78GptKCdwsZBEMr9ev33n9jNs
PUULfyKpqSwbDvfXIMjN5yA5MRgq+Yh6I7wnk6ONPgKNQk1lBWrHH0EA0JidvMYX
BIcoQ+8vhGtlEDxFRbhW8vO98ErCbuV90H9P1bfcvw5MYIsYM3HWaspMriU9r5Ww
dM+w1Q+LWV9i7tsH/bZsH4BT0gic24kKekaOA+vU/u3Npbd99p6F9CNCF0datqJH
cxyOqAdvTQD19DRZZkdtkHMKZzYzI5R05vSDhdaPLML2RGxGjB1XO6G5gg3NYR1w
3iCQKOtyaaDoZsn1aVkohIxIu18nj6QXl6sg6nk8K+ILqlKSqwR5GS1h7Uu+7Cvz
+2eDNptRx4+E4MDysue4MWxnToeMZba/xs68wgmGgJKJrEiK2ciCxrEkTHGhd8sX
nQXgplR866Yj6JlpkQb9Q5Zin/WKqSJNEsC5zl43r2bTvVaTXeY/GdESqcZZFRyN
rHLw7uw9IM3MzYworWVYpEc8m312rVP12YBRvEdGu2llahHr7IuED35/eIKfUNyj
zznrrHt8A6qpTXfEoXli1VelnwOR5OW60SkhK5CHQJNqALIesqpDOKoTTszS3HRx
hVBcNEwiWmLkrrCIsfQ3R/p9JWAQPwpf0AlLezLBmOn12pUlh7gs4IRsw/APYeR9
zaiJyCubWM6XFrwsaI5AyZDA+Kkxev7PYY1T3e4RmpCwCposVr10pUABor4Jh1jn
ibMCvoNvEPA8k+dK/nPEsXtGjyaFVFk3Gun1Avn7cdwDB6drwEaETBXEKK9QLDXT
ZL5ObfKosiVmjZp8HMAgCHPaTqsSiuMgWQhSb5DuOqOfaXVIf5llofMWkvhv58mW
6ZiHKeoHHvCiWcR2jgZk3sRFVEWR4Ki1fS1NSs/uCfwsYa+vmb4xJR1DaJt9G5Fb
yLKg9/Ueirhb/jGk9ZG4c3+DYBqP5EeudJyYsKot9Dw7EAVDr9rWZZAbzBqKpEaY
tmQTFknNOwQGBVMwu95Dh9sUUhxlR1Fhc9Bzq6Oa+UUnNiYgLMZvkonUlFFqGr+x
xUIk9GdptCyv9mT1C1Lg5DfnTNBFs77XOaDdUG7PigkA7LbmfmKa9yW3b8pQorc7
jGs5hAo5dSogrFPh1ZmnsnRBZROXPqGy2DEpTSyEJ5YASyQZT1N2BakoSXBaBeqe
ouaArIFo/IZZa3uo9prx//oY17r6F31rxvMU4glKY5ECmhE/Z1L8eBa8NSyca9dJ
GYLe2XO0VeqAYcUVnUlibmKcxidfgqczHgC/O12ovRvwjKPosibIFht60rZoLa/+
1QMcK5dAaZF6IIKNJEu2/1nK8aYFnpzEHNMbu38saQzs4K/8gIEWRd6uO2SMIg/3
gVHMjWv+zwHm4gFWT7Eg2C8itJjiczd34KLVKY677GzOabR0ko6NTOmBU32rHaFc
l+uGK8giTOrW93NmNo+7gLX7VBikYgIX1tIE4rOkmYwo0hayJntY2Z74PFSm/zgh
atIVLvEDUg+61SNkIE7cI5UYYXToWTSmaAQGBHZYf7Hs6kdlw4ewF7qELgJrg/21
PeIeUwWMkbCKPa5F2nA0HcYtui8HSy2/lRMV4BaOjjzq+Kpyf1u5qLvT4TUkVKru
ACNEilfLxN5ACe+6E5PFQqTMqd32oTvULtD+IOVF2ORFlwPTdAWnqNQOoIg484Js
F/ktwjLHYxbWoasnFvWkgBHmuOGykGv/j14Z+I77f5ryzDaulOGt1XsVhwpaLvEO
ekmqpfd0leKUJ+xeu1xhk/p/Tkuj1vZBp8BMO1zYxbWv34FLube9YOKh85LhQPnj
XIrevbQ7iL+CRIDuRv0WDg1gwOok1DQuBqSAbMd3YBS6at91TAB6WHA4kb9gqd9U
TiH92+ThbeIpOtZvUn/WkEpIN82w1YWQ/wPwZqEJeFocM55kUYVd1fTY92hX25nU
ObbF6KYpmbCTIzZCrvJ68rdxmUi3u5Jy/DF3RDmu/+h0sPKEJFcDlJb3dFTUt5KI
VdxbUbNwGE3jdQRiySSxdmQ66TkRVAIbADcchd7O9uiwUEAxerFSP682L299c5vA
e2DOivlqS0B8Jb7P2ZhvpS+sqJ83wr+czy1e6Mue8Ko8wmTRwrH5on4k4xNfugLm
hgWcF4xsin+LsgICt3hGQhkmq1FIVE2cKUN6VR2vPHWgOj689kMSn2rpfynmsN/0
ypGOFxRrSB188qXhO6mvvWMym/ggiHN6hMsq+bViSlm6MqPYj4jMdy/vaGD/ALo+
Eb+xshzzht48WdYIX7THxwCRste+Mh5dTWlDX/qbx2OjhxyYkvm0r/sedkg3b5bY
7dnpVOvrsMl3O0keZeUfB0iPhSaqhQVfOc/bo9+UfsaZXXn1q7BK6i+oz+7EuGS/
O9GyDVJ4Es1fVM+TgEF56WicrQyZYuBXTuv4kxl4HPBYaulveZv2/AYcfi6vEdGS
TiiCMK8ewwMtDgTmpl0W2Jq+6eytHQBn9geeZf3VPXhuB2W6sC2OEL7qi6JaEEJu
SALSXZmx9t3U9piAgRZ/oF1wtF3BOKJ9ST5yA6V33FImuyodzKYdmqxz1Ok5eC/P
ErLguVV7Uov1T4RUNtU7Ys/8QHs32vqxl9odxNtIn4CEnwR75TFS/Iwiot6L+Z5M
yyxW07LNE931X6kk3ncUJGtOfygROvwTkuEPteCjmrmBEeGX0Blb7znSwiPnqvv8
x/L/ZJuOT2N0vesut88QpMMgeEZ0KuPSJUXe3n3nvUGDc4f6zsrLYFTI4kH9SAUI
IvMUvoT3i5ztS1hV2f7sz3mf7UKnYyVj2w2BpskjX5EgFZPcj8UUR3nOdYcIt/g7
bu2bUq9i9RG3/jUuy1GGJ2enUVyaubw+3BiQ4ysO+B17/IRF64pZCSHwQzVQRyS+
p2mAAh4VhPvHQWICwSmJ58FT42RGA7/yZ+0WXaVfRBh7DLg/PRaYowDlARI7QAdZ
Ri/w5aVm0nm9dMoe9O6cjP8LLCqDxUU/nDG2ciJpa1jhvveQ5RuDWlPeN97E08Rq
7zIqau9xF4BRKZyn09UtLQVSCGxnxv1fh7aEOSVFdAd/eDUAvpKnqqN5ov0ibyRL
3FaXdrlK3XqLfEGz5QBKX9cEk7xjpOGefYNXrCnsI3QMB9kX2xliVQG3XizXcAGV
JtFTnnmdaJpiIirifOZCDB11zUdy5PUowL9OMhDU5ZB0DSxXqJ73ozofROwq9IEh
ZKq9E4uPTjNENZzzSX9zUWfFEmN9zQOhs9+7cClabJFBh4oKnC4QlOhOzEL6+SYr
tJAQKi+L+Fxl0o3fKQtGp/A/szUuJv087mcpy0Qp8xdZK6nTIXVRykT00980/0of
4LUlMU8h2p3XLluwvO4QBvPeyzWLK0pcYzf8Z+HNHAt/6yoCPq2ry3zPBUd5+AyF
cMpUoExsbZUbR6NEh0oA7RdG/A0POayNoDibLr0xeZ7yYuYEMG5+USkl+WmtzKvj
l0leEl7nEEBKxP2uHsvz2PsgZW4y7a3xe8PZr5L4PS6ehGNC4FMllYUQia0qd1AT
CNm1Lgb3ZZD2SrTkYbbMD5vbeBKgulDLpKd6IXxztXMQbAOxDR1lXGxQADNuzOoJ
w2pJuCzpvxOH2A5c9x4HE5yBtqksbiVOsT9ZocLXSFOzHBelBCQ+YfLHjK6NEFgL
nUVbA6nWU/7ctzxfk7YORW6KcSw8YpNVWmxB+NqltAz4romMNTACq7On7Pvafc00
pfUWixNRRXtfu219rIPOhSL1wnxI232UoTrhePY78gOPckQ/jL9ri8R0oSrfI+86
8t7IoBTSA4VLQ6G7eWKXxm78MWPfAXu8Eml3sDI2avc58TVdE2eWw3QyhtteVNcB
TAfeIPNkZHrVQ7C8d+iGPqs/eMs+y2BOJJhhPb/cvM/0Z4cO3cplGKzo0Fod2/1c
M8wY0Aefsh7copTXXk4y5WEt2EL68tJBlDmmrfcjlFtyMFXddFY2ugHiGhMC09Fx
g9ZZaSKcB1BZlHBQuHdQ91BrPZ7FgQVgi8w+y4YSyjfJ+0CkjnHeFl82sqIwaX9g
FgOQj9kLAYSHiLvqiE/rV/HKDh/zNGn0QqfhPTjBqsiXAbA6Gh/N0EiiUu6ZHOgK
btXXEh6sM5hjuS8KUQcHjKqmhQsTSH5zS3BACxNVI0u+6v7HGT2Q3nAF3Bo2yq0t
XlmZ0BZmtWhwg191H5DutuIPJtibk733hHXaQZCTRvZ3Q5pnoSCxOy7UNH+T7h9a
T0fkelNemXV9Hb+Vi8GpfqRRDykIdLsCP7tNYGWkRJgNIR8MbsKYYikIbJSH0Vjv
bgKAjD0hTuIrO5GtGlIzS/oShPn7JaWPjKBKii5k6cJ5Gpdwk8YF+pbsW5mSbuJQ
lr7SaPBXzlYhRIJnUPrToA8EtRPidaYF9jWq6UKkaO7s6i6x4o/gUjCufsBuM4r6
hgvSuk7SP6D23/rC3c8Tzshh6LB22/5ikLvDCEOMDivWEkN+maphGBad1Je40ywX
jD85kXNkchf8oL53CtYNJYYj2oWC93n+oYvXPJuZTJZfBgGYk7KNWaj8Ktt1rpyQ
0TMBzoIAx4vHP8DzPbmM+dvKDz/hdhkKTgYDcCk/xiBwhIZKyglMJ578XzUAoINr
glLk80gvb7645WJ+noGPRrNw0k15+rc//LkF7DOXEfO1e+jor0+nd06Z6MrCQNfn
SA+lSc9VtRsKi0ywK1XVJ5a/04VLn1OBwkNRbdEkLJkVvgW7X4ZyCPkKUgTCmO5x
9kwMxdC4i+UgDpdYMtCDKxOkMJemXW1ua9JjRBnvLTxFeEEv37PaT2X0bibiE8Ph
KYVCQoBIyzzxUbdCRBq0xS+uMVsR6Fy+dzLOJr9LC3dS+C6/2Tq8HVizW66/Ya6/
5wZ7Vma+fQXHWmKu581YopAQk40ymZ6hU4VDy8pFVhClEalk/LrdzOEX5tXsna+E
osnt468GN29NH+LBsayNI0g5LP2iQT3B/Jjll64GXfE0avESAg7dkfCd92PxkeSp
dDbcAgoCZczTk6Lf1qH0lSilpjNImmS1mtpQQ3C5jCF0aFRuX8otacfd3JhR79Vh
1ABn8qQUWx+0TiJhSGMdcFEMbrEy99N1qMYmVfx7Nvwo0RLjl4fr5XiXD3UmOMvU
If4alSBdkmJ6YJLRm3Sa3ejEajjdy+eJWvqkbR+d8qRWJAB3k+SSzCNSukGavBWz
lvxy01b0JBVkUDiROs0Pp6Vjh9viQos03H8EqZY9o+4w+23/o61Ft/X+zvFCrlsa
Y7wRdXlxKIkQpg+0PCVD9bLqZZcNWPhmblbzpUNprnJ/IYSJNUMzE2LNRN7ywSxW
Bnh1tlOZJbyO1Fan7YWCjEC2pZvOaH9XUvbkhFDgCavSsmWOrO1iPZT68oSthuJE
aEs5N+tYT6WLq015IfbuLWh7HYd0xlV0H6aA1K5XWieZ2wiujTKIdOUj815RqyQ9
njw05Y65NZyzvCIVb9eyjnoB8hitefpd5j09o2zR8ajVdaLfMluMPBgphU4oROeR
uPCNK+j0fUcnFwDZA/WFFXqyrrfOUabkdk2IB9lgK63WqMxUxadplustM8YFZ34J
EijCy+LzSiUK2nzBKg1Ydau6utI3TTh6lInstjROIRa88UhHlcz18L9IGEhWVufi
Qd7b/ymKKcZ/RrDPUSegJ6UW/OgZG+iXYDDg9y86MNLZnRuLOWKX0k3NxgJQQK9V
LbM/24gS+CN2GFIcPRM2mqf34lEMpGz2RmTmPGqA09o2HPqrZAUStUT/PrkMfbuA
0l0Y4WFKo7EOn79Ha4Y235J/iwiVUJ1ZLRuIkcfhqsbq+POirKKObNT58eV9FAlM
lN/fvjjmbi69rIQ2Q8eMHTRnAk3zKqmJJ75Pfd/7kWkSdYVNT+jdOOGaeffTqTGB
9Y0w++Xk2plQ414WELVPCKOElQD3aHe4Bs96mHErb6zWmwtB+/9gjsHeMl2VMRcK
Yw81qi6yCTMGbAeelly5NwOBag5kBeYDZ4PD/4d3oyiL/4lN4wklBSwtoYLInNEr
n47eHhF3jAJsXZcc0zy4o7jgNQ/xeukhH1mAFw25RLZqxQymoMzHq3jEu7AAx8eU
c/vSYIUNiSSSci/4whZQcpUxX+7vbYBbvyf05FCfOCUyv/UVAjXCnUbn+82cM5yu
fGuYVohA0NqT+IBefeuuX0XIKYXuRdihMfejaIDjnUGoLptRQlbwcgVAe0sFEdaL
fQ6s+SU/5gK9Z2BDVgJqYDqy69meZJ1Cyih33NyNYTFBCuNeaUEUsktlLgWLHtAu
9/empJNiHtdstRzw1JEbNG7ue9eo3FC8fdB0y5RdaEG4jwk/mhAQJeRmAvZBToKW
0S2UXZ9+qQ6uyXBQxQ66iOylKOuXLuSfD0NrYVCsGofPz3s3nPTB7pA3eb7cEHbZ
lBweqcU30CGJ9ZawpTFazT1evKldxuKrYlESdfQ4IHAmCjBZ/QCENOB9drSVykJi
0UU/QxMXt3YZ02x+E+fpoBWHPr8t+d+Nok33+jfFp+hT90tKzYAVxEqSsntiCQPJ
cNUlFx53WLCQzagFFSyb1jmekD39wnObiA9S1/IfFPTjPF3/ISjvgvq90ilUdIIt
AXDIX6jek74Ebu305hJCr9z1mZ8XUCPy+xNVvYt/eWQ8jCnVC6kwUXssJcPmtzdl
wRQtDnxAanPKOJ3XfnhizuInVcQMNWAk4JstcJFt90+80bI8QDZWZQ0aDgXN9ezS
G9z/e5enKVy5+A+pl8poXn1rwB1YNMoHXuX1hXDIaopIeDFv5uJLgFvoCK4+g9wW
BWu4T1MyNFqUTcHLc4vBlJesrRSz5nB0x0SskT7K/i+xMjx0yqHBbmfQ6xkJPj4e
DX02GJ3+Oy1ofvFb1L2OKlWblevx2V7q7fWT5fAJuCFMqqGKHidRh5iE4OFc6C7f
vpH+gws5hNPuTAAu/4RQmHkLlhOWPm5zCBoYWYDP0DG7nBaqrC1CxaosHkCsFRim
B89P1w/lLUheTK7y/zLiuetAPnIFEwmuT9JJ4uqLwnjaOA23rhi8id/IkxxpQcdF
Wc/mnYuBnHG/cObU0Wa5KCRIpHl9DRn0Bn/GfIKXuqlySZX5sa+j3Lx0xYLW5LoW
TVrrIvDdC/ZpBEcwt3rLh2wFeMURXwfRStg0l1H117A9BYBzChzXuSN0s64n2/jj
iCCE3nwr4qX6zVAwvVcHA576VRDxOxNqvZGoMuMPVjzY+D3AjVvM+pG77X46Ar6L
byzUnvloHtdvQCL1+5Ahqagj7p/YsxvNI6s2SEsccuavKF7hRKCCTwshX2Zhqxd+
HwEdIoPlJ/eq4cHRYiIqIBnAw48sXidXjO2vYBZAprSNzFGPICBeTl6YWyDA80Xx
BctQtf+NF2L0kxMOuC4sSy/nP012mmFrx3cB6YJS6/owEHEqFAJr/SzzkZrMQQ1H
BoLaiS9MjGTc5+gLzj+mPlEez8Vk03SyLf/tTNeCr08VDnhc8h0O0IzYZI5UUwCc
Q/GIj5v7VO09tKXyMdwjAGetMrHSHPUkcpIplOINQPzXQgJ3AsQDZ6JHVGzdnD7r
D1fjQ0XF5IiQlXFqFiIiB3RGP+EAPcr9i3UumFJHJFzq2TwihdhtRmd3MiPTQkhq
argtCIw+GyDAxika0uKSkhx9/DovJmZtUJfphj9wwRU9CxzbipwcglBdrKJvO+3g
ttf8XuyuEaKuYbJrXMrMOdvYwsAeIO9Kjx36pjPXObsSIsykKEOQclR37jDIFWKm
7nc/urnfLCCFD9XvrLQ5grtCmR6ckeZIFePALtj30AA22Wn06RI8++mCuma/uYNK
udj0c5ZCp/L/35AmGfxDujAgnSYgSnEJqnU1hbZSk0xXkU2vjJ4Jrnfvn8KqfRp6
H4qn0jim4xFX9sGX9o7m3WdqcBmFKbGgdWQvsy4qaW6MPnMdERiaXdIWBzjDPHlP
/mjIsRLwRxa+0vPtSJshwD+v4U8jJ6bVRUrIVwV0lF4dqLfEFN3dE2Glvdlo7v4Y
Wr7Grgx3w9+90TqIPK0qPbZmfBqLuzUapKkfxxTDbPSskCNHZ96CJdVSyQCim7Lw
qpcS4X4yXJ+C7nG+1NQxVeKQDXfjSDxS6YtdmXgubr3u8Hh9qMzAyVTNXBlc8SWr
vVwHMM1vK/jeGDzGGNh5as8bY6gVU1gD1ifU6tDZQmqNC4Co4E2gMORZVC012rLM
34DbxAGdkz/hokPS95qe1dxoPfaab+ei24SvsYAn7UoMl7LUBrUIMDcCOAl3d+vp
18KCLWcN+5ykIhPh5XyqAtDHzIRRz3I6iNh7xEKGdN9Ueu42JiV9RH1ej81kCCHW
+u0PTDhtyOMNmfG5qbR132quTQ+OoUzZp693bQn2PcFNdBbrVwB5BEfAS4msMn7S
hV34Y32wE/5w60SX6oBMyCTdm/PVSISYcyzPrjtzYEcqZe11zCYDBCjFyN665iAF
U4C47tFDYVkMLMsG4EiLlEYsHM+1vhbCTWr3McbbOCQOwHZotYyBz7ZUgdxZfz6e
rQj0m1R6f8Z9+X6AGtUoRj+XvMQ9sKnud7bt8S19CsV2+bLlhcZ5fkL78y3+AYRz
a2TUoYZHU8idW/Vs8DZMhefPE/V3RxhHPDFlPtPOlOw0S24NyAX5twF2FIlbvLkv
dxLot2Cx56u1xE2sBti84HzK5/j0WCeOyZI+kOQqxT2R6vUVpTa6gKBL//c3+065
Goy4wRebUXYKuqEvv119ps2oAeKhrneISXuS0FGk7pZyIpQKc8P8J8Cs2dTWPUNp
LtOPs3zUtOBpbc3ImK57gshTUHTouKD3eXSAvSXCFJt+5VbO+Q0fr0Re8EBcu7zC
geCPoumNL76RiEAmJZESVfQzNEk09rAGRWZV28hX3FsB7TYKlSMeB4G9yXiNtG/g
8ZrvxljD/KHQcrlEQfQ+2ufBdcq9mfkHDmJSKf/Ci7U0pQx3gLS4oXN2P4zxhQl0
N5NEDxaR4K0O6OBQKVxxh7tWO4C19Q4lBVIsmTSQfKIt1dkmuYDNSWjxBS+VZY1+
T3UK4IbTiaZw/UiuelWYl0m0yX5KkJS72Wa34tQPkFwOsz08UHIX01pDJtx1NC0h
++Wb6a57xNfJP+n8fbYTe8FVaWQulPqzcj0cB71vz8ydoltzq4TJsgUYkCgHxo+5
ub8G863YA1ql9Q8ZNmRw7BGVlV6gi115ICX28Sek/5nbCxR3dVT8qDXeNJRHCcyk
kj6aeNWFWnCuZUufzWV9zD0MDnM2bcHvoPkmUDkaPjtXU14bbBnvokGaytOvsLXd
7hkEduKdU89ifzyuVwOqhx2q6zEuoVfl8U7Wg46usSbKSWOZlaj736aprs2cDnHb
lmA2e3xM6db/paMlgi+1x9/agEFFrV09z6XwY1vahdbrUeVVdubFZfRcI+WtEGaY
uPUwt67j5IIEmn+Giov2pTt+XSS3494EfpxHStKxGYGQHwyA+g43NxCq+8TGI+ma
woF7+7Pdecw17wsb6Wljr45NueR0sfdiqua46d2IvW+aOFkrPe3O/6MYezv5ZKOl
267Q1z9b7qqTLw2QsYyK4Ob9s3hgWunfyoyPMV+7GPZ1CxSLp0TApO/dU4waYcXW
4v1NvRQal7/9U3cPbivTiJfqctUFjSsd3Dyu+vmiDNin+0BD3pqgYhYZCWAiIAfb
UWPn7gMeBZLs63kxsVr9hlTLGdTuIOIhTNRTYjwN1dHy7hlaE5HPhLA8c4KBbv+j
kCg6GmU2Cx37KMCkL9s0o+foL/CP/6VtcIBMFSmjJJyydCKd7hXNwJ4E7xKBdZrO
sq83Ul0y9CwetT2NH6+TiTmJl5PmIHtpsvxQe2om8eAgk4m/fsLhoaixTBAlCXu8
4a7Yqk+5tnTxxkk51GbICRJ8/G3+GRqXiBl+s9TDHTwzfnwJrlbKRKl9Tn0LvqT0
slyyn8CTa9E16fsmI5EKvs/yJ8LM4CsE7GDSnZeTX5iuMGy4T7n38exMb/LdgwzB
fiqGC4LGZdD/377md04pLXwg3slJd51ggrg6htaDOYg+31OcjuxqobgjaHC/AJsE
gDgqEvhc5nIZCAKPxGUfQkyOSDWdi4d1r7sliDcUmvWHzNzeUUnECUeXZd2XPtmO
tkCDYFOYzfR9Koi+ajL6lVWFHdBogG19elQ7bNzDMUMZ3KmZ5y+t9XWWm3fGmPIz
LOm1uA06pfVF6UXhpduCgci9t0HwDX9hEWnvoSefs/3+49hTcaCPFY7z75vnTgh6
AZDCkp8kmUbKRnjrnzb2N0HvdvuEY9BmbSKA3cRZvIu848fkykaXNOwzDAbAxTD/
GHtFA14J9s8bQ4jMiBbzpRIxVmQqGw1vg351J8nAKGesZcs0BN3EHOZ6ze1WhnCC
BdxW0rAdNIf0XmcqsuXUCMxqUe4OCMmw7NAyAROmAz83VXogNJzzT5QQ+wQUGoCO
KqhuABSq6JX8LoSgNSS46vhtKpZ6R49V0SXwSL95lrISBwXTp0/X727vE42vxBrc
KSLHJFIPc1RqL9VeHGFIZx2JMxCgS8Aw5MzfrmQQcRnpDAeJuDsWesvFf+IFeKpI
7d254hIwyoDiBc8fcLc4SdWd0oApkIBmSQ9ZxQ7pAY18z9B/y2pf978f7SjR4UUi
TRL1thPl0GcIJ4YNQTDF/Q1SNNDMHFmn7AcB9EkgqoHZEvODdFyes+ZshWDkR8vf
W2fp9UpP9pLMt0beOSBjM4nG/I5g+nysaF9rJz0Q1eCCxO0V7PfyBAgSL70sJIZc
xL1fFENu6L1T95cALHgIE3bUGfp+79hf+r3BQaQ8SFE6uJqrwfavc8BY5m0Y/ldJ
qwPxXn98flg30kxHnO83XVcpkW7K2xfXvUKpQpIpnwIoWffRVryp1QXRQZ4k2gx7
sajCeLhERQhVsbg0/1CmhB6L9/VwfhbjB6Ny8KfHr6wYOq9vrpX9iXbqaQDxyJZa
IgVZldINQsEzy4PLsFALRMaP9cUD+gm8ad75Sq09l9o0cDslQ+zPmID7wyOeogM4
5YaBSma+PE6atF1xj3VIY3Uw1E5I9+i7AGwVd17W4Hti/jxO57lgupLIcfqL6TBT
RnmMMkYyY97rzxwLGLsY1tcNEfdxPq7ddxExUgUZGvKF1CvgEJbkRhHliUP634Or
m0rsCCk2kuqkyo3HIVn3OcjaNjVjgKPQOlRal8FgcdjCegKRdfK10wtIsTlilAKg
hpKQS+objn7nBWIg6ZfOkDNGfyTnBnMl0Hh/fy8FAVPPE7gkFSvCW7J5f229xP4G
QaB4aCWEEH235X+yL0n9hA/nmFE4PrLBqcL6+hXcKqO8om26IaEhIMmD15gQdEKi
WhoZ95hYGgv9jTURd2SRHJsjhICpqX80xya0b2unHVKheoxmTYV4ODOvGUvdv5v1
6nES8jGUU6sjSYShASI9zZyHW2/CpYXy47KuE1FofpEUmwAtGfWg1hiszu2ukeEh
04B4TN12BSEW8/87Eb0lrQ/uegnGk8gwCpFES9IlEZVcyYdWIr9kB5oG8AA6Rm1j
juPPCHTAdVjCdtE/yEY9QpMK/MlU2Fd2PinvIyfPOKzPP/xjIUF8CWEBpNf/5Dmk
kScWWLW8SmZo3EskdRqwFNgk9WFHj0XUcz2/p4E18FXBCnKRlNSsLy/sng9jzTF5
c0oVzbAWASPGeH9Mof6bwNyhzZioHzsHghCe5bDjN6s8QIQ+Fsp+oQaQ9hgEBMHw
ab4zAnb3Gun2T55/eIU3yv1N9HV0YFoxgmqNdhlbpYSwaWqep0+TViSFNQqdsea2
I+ZttFSFTEyvHiiizJFR5Y6XxMH8N/9t9j65taknDHffKbXUzRSaFy/tDK59vqBu
JiAgRJ2sy1vEQ5I25yOUPBF8gQezDQiXWH2kmAv029HVbC/+y067LI/Awe1FGPJX
1n7UUIcKWTZbNXJNUGHWXG+9hwa1eENdinB2q+29tSHJp1BDsaXEN31dfBXyuIEn
Iw+ltSc/4rbTrva9kiSHLZmd2t0SpDidBkOVGUlL3Xt2UiBG0sBR9wxZl2x24l+r
Pv8KaC/xEQBATuq+MFUUSlS9Y5dO4g3ffnxqmXmO/WJ+rSyU9dab6VF1nM3ieizE
CB5fctvHjmqdp/U//VpG0u0AAw52QOK2Fx4ZjhYjU1rvxVkQVXDvev+i+AFbbP1i
zEcu44ZDHMSgqNUHHU/nkp8QoAtyOSnpnWamHpJRaZUEBW5C3VebFKZmVl2BU++8
Mk1Eu8ZQ+5vfvJdOEdweQvadPeaxDra4W2ZsP2Frb41y+IPXAToTkAd15QcvXOh5
v+ZgOcdG3WOMUW48N/9ykSISi4G+AOQNoqJqNeUzysYHp2Pr09NHtNprpqCvtTqK
ks6MpXVnwWVYN9veOR2sBMPIS/RvCRHIabcRytm+lK8WCeRRpO4mrxtpNNDjuU3J
O9/i2IV7lvf9Q30zas9qT8Y9ArLD1pXAxzC+sOIIv+iIc0/ML94kh6AxC7+aPLTy
0c+g50jUSz0MzfWg6objjCMFos9VEZ4AA0HWDUSiq6b74SZbalTZPijAjTpG1XDX
auxHCGU7KaKs3+NhYBLbwanPzAGoM//fU+rvfpiuWl1XZ2QJRAcw9MXymGrAzGzR
p3PDLFk84PQGdvBSEQJJ2YbU31ktlD1JLX6KDpsZu0/OC7/Bd3IiBzBQhty+N/p4
f45HZMetDv4geE1NL8QGZYYiimF0phzStbZ+XKD/Vi4a56ob01ududqh8Y5eAkqb
VV0RVmiHAAo64H0CDJn9weoe35zDzJVdQNQl1+vA1va6ek0gvdzaEc6XnYvtzmgj
STsB8M2p3NGYF0jEuScPWPpJeqBxABqKaUqWTooAgnR4+VIau6muDCCCK1Q0hKai
nVLs4O5+BRR8vCS5HFwWwRMWfUgloeIi/M49DOHMj0xdeLpDfBCubCJuV/VZtTda
kCn2RrROk2yYTcmpNb9NAOEAW0KbO1A0fBK8TGqZ/eHWkpq+3WW0rZeK16U9wH3h
5T2tWAoiLla7li8NAOLA7JdLL42F2CcBTBV+K74vPFQOShlU+mC7BoAf6SCM7nLF
WDi416ValJo17flOtEAjd3d7PkcDEWs3BIZgDcV35yMZQZJu/7Zr+6MsQjMKrDEs
xLG9C0nig2CgnQwyDTbEZKqzmvcRV1iF3E9qfb4suEQ8duLTXjH5HaXt8jgs7VSY
9j3YiXXVfOnmxN/QgZw+BN5No7DmPr9LngT+cVM92UCrJSzHqV6snTHpqOJSvEgs
o86WAmyHqwDZGa7Ii46ASimIYNNrQPhmZUGXXA6XQ9E2/s39bQzFA5mn+7uu8Hnv
oaC1kzhYfnlBgBRn2TAoHWYbfMNzcR4AapUFD3rW0dyatd6+RbFs1MxH2yIyXapT
TeXK5TrLWBl0bCE5xqTHi4sQodotDjzoffPPEtrkmf697YYz1fgsldZ/fXHa2e4+
juBpkmayBVeWoB+YgkaKV4Obds2+COzlcD08pFn30XDiMxFQ0gneF5ZDcL4DVQwX
L3pXJbGtQfGtrtM6D11JyYKwz9ApioS1iT9afjgfnBDPq2T8HcWqKXLpNiwzStRq
MvqZXVbUEPNo+mcaZurPhnSc9KCkehfYaIzOc+VOdf5JZj7cZFRQqVqpyxeHAIZQ
MouKOKcdhJUf5slHUlB3sDeTonp0fQ3rlqiFow862ZEqrFZYJIJzQh1TcNHpT0d5
2F3GoufTg3e1TLxE26ef+cniZ4Rc0pYGYYdB9p1Ny7tRmuQdZhn0y+/wmyJQUU1n
torjJI54jWTBzYpSrQadbuTG8MaRZi9DHz3Y60eEfwR4q/4OuD8nFww6PZNPe2cW
CPsYL2wuakv3l8v7E2+wWkIuAPnzImXjldSNI9nQElPGt5Wnu4ZIPsrQpsKiuH6d
GGq9FVylq9EMO7/JLYk/ZRpK93I/fB+Zx4B5Ibi3hjWXshDEH1j/NbGf9mDB9lot
xK5jIxf69FMhqaTecTlrPq18eNE8QuRrtYv1qwX8VlifrqBYtMmkfJU3dM6rvtXA
DrshyeMVTHLh5bq4nu5XOFK2raILbA6az7V7FIneRb8gws2QHy6iQ7ER0T0f249S
4r66lTBApfLDOnhwlXG5rcRwju3w3acE7RjqnAEjDDXD6gJfa1SNOV6CFtoEK/VQ
OZe+edzk1p5Yr0m31K0eOkIeCpLVvL9EQBAmXSjZVU/8odrjc3kJBqt6mbI2z1Jq
c0qTIfhhOxIxIGXpy6gBd49lOf1rBJBpMowrY5btdJOSfJYsf/aHswedTRnZuK2u
dVHFRcjpwci646JrOceA94Ayqn4aMy8efjc7N3cBI6CQyExeINdUQtgcAeH/MLv8
a2j4s8E5a+/VY4D+HxQe1edNJurAxaqaXDUwS9O9H3mXeheKbOSIXYvNbv5HWCMZ
lIqRRpnnQ4IrsDaGey0zu3J9YkL+w+FMUoRRMGXkL2+Th0zOhJLWlV3YS/uvmqAD
DmWM801RgW8kvPyFHPC68zj+m03imUAL9ixcmit2rcCFRzciKCI37hfJ3mWEcK34
mGJqRKtemtW0wfH13XKZ7oQYWpp4Lap1ESwvhDSwsjFQ49fOFuW19mrPIw58CyGK
FQ4jUHq0ZLh7gxWWuJZkaHWSvedR9i+buz6Wlp/G8CqENvH4HO4K40oJHtbIpZbF
zEePVsl5A0vtYYFea2hL7bT0aFBILY/Qm/ICELfnBkuLT/O3LbLPBk9zKfmpw33+
SJtNN2tRp3iMC5RsVfvdekLaDTJCbEezFdN7+D1A+KM9wXBDIwWbHH8GJjx6xkXn
zoPaqc9NWDDgSHMLZ1H9vlV+rwKTMHnLBLwKC/bhtJpIWkJj07S5aEq+ZCQtdnG0
TzdS747EWlapw0cUtiiVvrVXM9CPAI4NQV3pjOf0O9fso+n+p98PqSHv5GYnwgZO
oUbvW5QNOwRylEIUxIUCr87SA5vfXU5BbIkTMti9jn0mw4Tog7SWCNu8PbZndyqZ
vtI50Nr9B/EvDWl4KupqFBba9YCHkru1VWMzZjPiBj4vLe9V/Xv7NNYOufKNcK+x
a0jDwXThGqPrH4fcgFzDl/bdlyX88ilHoUBe7nzTlWcSxm+6ZRfb/Fwl8FybKKza
Xx0LqfcwcaLCYUQMyMfQ/EG2iYPQnsWvil89/CcPSh5YU+G89uSc1ZiyTyfKLrHO
BUJOApg6wH39LewAvCI+7oKke3WUax7/6yxbzOumdy7GHHYPNo3B3cqtczEpr301
c++wyZACZfqIgxWgKVinq47YDd7Ss7e5d3iaBwa1741mOQrxYBZiEYQf73g8V+JG
5Pk4qsUeFfIsEqVWytqubA7CRcVbW3vuCmVVN+5Yprswmudh6YfVMeQfc7fW3HW+
nxBhmxFiQd95HHSdWIahPJzon/JpQaMCfXS8PKCG+JKDLmpggIMj3TkEqlm3wDlc
1ENKgc7fPRaCYHuAnRwv9poFxQ3e7nPrLbqhT/xkRTpQ5nyVZcwNB27euvvJfewr
b3XQqSHYpc9XAwW8GGhPE8OX5wrdVSh47OkgxOZqOS5wTw9lHCel+iM3cjVxookm
rAd3Q0ia+oV0p9uP7Mo9F+4HRro3u0LvBfUlBonQ31mjPkzDwKvNjSUrjjjHz8nD
VPHrHat67CS9EvryJsgB3p7ARM+kW6iIELcwmor1WMpPjhiX/4Bx5zoVmMnIUWrS
qR7e8EmOi8Vw0heTlVR/KgzV21BhueQSqejkrsLNNnttqj8zNzCBc4ysTCiqBp+U
6jGtAPzGs0600OjTi4isTn3lHscEHJd56DzTpFfJ14x1jcO7NFkCkhqw6hoM+O+X
1a5R4zJD7c8el58pp5q8gH7USA/REV+nQXDVDhYmIyMIvso6Zy+SE84yKoDJUpta
Qtmrf3KwhHG4dqWQqtqjTfrpK7XakF7lpDitWWviuneNrS7hXSveMCPmRC9nk9+V
+H7JaeG7jv8B0BtKS4oCXZkQT6/c+he/gi0RxR8M6ar3ifAvrZIn0rH7acoXjs+U
jQpDjpL194HaS6cYFCDfLg==
`pragma protect end_protected

`endif // `ifndef _VFLIB_SV_


